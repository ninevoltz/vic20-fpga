-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.Vcomponents.all;

entity SARGON_ROM is
  port (
    CLK  : in  std_logic;
    ENA  : in  std_logic;
    ADDR : in  std_logic_vector(12 downto 0);
    DATA : out std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SARGON_ROM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'    => result(i*4+3 downto i*4) := x"0";
        when '1'    => result(i*4+3 downto i*4) := x"1";
        when '2'    => result(i*4+3 downto i*4) := x"2";
        when '3'    => result(i*4+3 downto i*4) := x"3";
        when '4'    => result(i*4+3 downto i*4) := x"4";
        when '5'    => result(i*4+3 downto i*4) := x"5";
        when '6'    => result(i*4+3 downto i*4) := x"6";
        when '7'    => result(i*4+3 downto i*4) := x"7";
        when '8'    => result(i*4+3 downto i*4) := x"8";
        when '9'    => result(i*4+3 downto i*4) := x"9";
        when 'A'    => result(i*4+3 downto i*4) := x"A";
        when 'B'    => result(i*4+3 downto i*4) := x"B";
        when 'C'    => result(i*4+3 downto i*4) := x"C";
        when 'D'    => result(i*4+3 downto i*4) := x"D";
        when 'E'    => result(i*4+3 downto i*4) := x"E";
        when 'F'    => result(i*4+3 downto i*4) := x"F";
        when others => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO   : out std_logic_vector (1 downto 0);
      ADDR : in  std_logic_vector (12 downto 0);
      CLK  : in  std_logic;
      DI   : in  std_logic_vector (1 downto 0);
      EN   : in  std_logic;
      SSR  : in  std_logic;
      WE   : in  std_logic
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
    rom_addr              <= (others => '0');
    rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D30F57D10B90222A8593546710D5D5111374382D2783285D611308E04E35B113";
    attribute INIT_01 of inst : label is "8723080240C589001404005C189856330D08C50822E621888618232085610881";
    attribute INIT_02 of inst : label is "50720EA0C812023839539161886C8B9C01320C5816C480385E0441C3304334D1";
    attribute INIT_03 of inst : label is "B290814505C112E6B81145AE1084804DC732C6168D5517175453454535424248";
    attribute INIT_04 of inst : label is "51851D2010A04838112D2CCD26D2331683168315831780A2475DC74D550002DC";
    attribute INIT_05 of inst : label is "75DC74D20A098B6D8A4E1461474554D51810D55B55544D55A8DD920A22467578";
    attribute INIT_06 of inst : label is "A3740111374A4F2D119DD062F2B7CA11D120B289248D75071DC72F189D571D04";
    attribute INIT_07 of inst : label is "D113308A075DC6CD0A53496103C90CBC4C3477001BC94C2D5D15469A970550F0";
    attribute INIT_08 of inst : label is "36C00064703B04E3115700B00621456D1D534745542055BCD1D5F34744147C19";
    attribute INIT_09 of inst : label is "64447414066881B974466574110D1D14F07744435747143CD076314C121891E9";
    attribute INIT_0A of inst : label is "00FD550000DFD0FFFF934E934E934E934E937E933900300DD5D019D1D5140574";
    attribute INIT_0B of inst : label is "00FFFF0000FFD40000FDFF00007FF40000FD5F0000FFFD0000FFFF0000FFF000";
    attribute INIT_0C of inst : label is "FD57FDFFFF555FFFFFFFCFFFFFFD55FFFFDFDB2A8A2A282AAA0A080000FDF500";
    attribute INIT_0D of inst : label is "FF2AAA0AA8FFFFFDF5FFFFFFFFFFFFFFD6FFFFFDFFFFFF7FF45FFFFD5FFFFFFF";
    attribute INIT_0E of inst : label is "8370DC370DC22F881C53406F90C064064ADA741C3DADD00000097D2E7808083F";
    attribute INIT_0F of inst : label is "5E42F3F891457507155554D564F6354D6541C89066550E931506F901C53422F8";
    attribute INIT_10 of inst : label is "10455549A09961B49C8B3C062640502C1909C82CF275273011CB15DC24CC1955";
    attribute INIT_11 of inst : label is "654E1402003451C03C22944544CDA80403770DC22445114F4C6D046907984918";
    attribute INIT_12 of inst : label is "8C9B170732880024919718E3DD718243164023C4057221130F4142E2C2303108";
    attribute INIT_13 of inst : label is "0084E24CD601840D1134744A30344362004414005D148401D04845987038461C";
    attribute INIT_14 of inst : label is "6349802B0546444941054281104044A18408242164E04459045C0615A2C98D26";
    attribute INIT_15 of inst : label is "2411805D81E3D9D04814D14D134455144DC40A227780D58A9E15D4D4160398B2";
    attribute INIT_16 of inst : label is "B5D6B594D8585DC4C4609320931D144050840E919F040E31DB7440289DCD1214";
    attribute INIT_17 of inst : label is "920A0DA0C90100C50C20E6F10D14A10088D104610342220D19502B7537171771";
    attribute INIT_18 of inst : label is "2F358038F374E2089274141126226138F047748C3A8B249E926A58426408D042";
    attribute INIT_19 of inst : label is "448330B91C460406D44890891210183C193003510A00289D0702930BA28C5BC1";
    attribute INIT_1A of inst : label is "4D44935E71C6D1A772E69E208321891DDC8820E2142188308C85086005458005";
    attribute INIT_1B of inst : label is "80C0D3062892536050A05130090453634BDB71F318590F490E450F6D0E690511";
    attribute INIT_1C of inst : label is "63760B209224C20C932434402ECD095899015677373609963979ED13330751F5";
    attribute INIT_1D of inst : label is "433B9C5DD9C9CDC279BC17D11377459C24C90910A45D248A04044DC5C5933343";
    attribute INIT_1E of inst : label is "112301559DEC59252CA0E1367099490749B4D5D99CE3B49C125A248D1D990354";
    attribute INIT_1F of inst : label is "5E23478CD14D45488D505189088554515DDCD08410B8147036099628979E99D1";
    attribute INIT_20 of inst : label is "2C72274442ECD265891E5E7B44CC22C1D47D6233B885DD4D4279A77470257841";
    attribute INIT_21 of inst : label is "C90192321248CD5E74679BB2564CD9868D1050912A2446165542663504445353";
    attribute INIT_22 of inst : label is "5D42088E70604D92246717514716148451412314536711416434891905C19C15";
    attribute INIT_23 of inst : label is "146227794DDE7144D9CDD249C5DE40779298D8A3395298D0DD27B277496DF47D";
    attribute INIT_24 of inst : label is "1A194102AE451889DE5377905CD04DD24D8D7374909D25377981DE7A44D98A39";
    attribute INIT_25 of inst : label is "39242EC1D421823910873755AAD40C18D6520928D5DAE062826DDE7911D8B595";
    attribute INIT_26 of inst : label is "8D4A89A4906054585DE0756516643855D90D9917538A8DCA4746544F6DD24881";
    attribute INIT_27 of inst : label is "763552757304D204108E72404D960CC948588180803D034B5AA2351916B0D6A8";
    attribute INIT_28 of inst : label is "D124491044D535234D0664914D48D3948C3354424284D1356161241509011D13";
    attribute INIT_29 of inst : label is "56088961540145027174959E1DD959137412A154A85540912647655745491344";
    attribute INIT_2A of inst : label is "2350440191949852336466143409459315485C11008114D0112246417271A929";
    attribute INIT_2B of inst : label is "33748DC905923042706409419305481C50190050646606409499325489CD022C";
    attribute INIT_2C of inst : label is "01C9011301105434264CCD49185DD20414336D295115D99AA9005177264094D9";
    attribute INIT_2D of inst : label is "405706245250749330417014D1C941301414DD36362624054140404142463617";
    attribute INIT_2E of inst : label is "14890890585890890127490D27490D055D105D26933240501933053474061462";
    attribute INIT_2F of inst : label is "C945D274492D1D518C5247491D2DD404454D1491A52C410124964514D4905535";
    attribute INIT_30 of inst : label is "5152444984927340417413264537349125457143449F4927D2506D0F4755CA0C";
    attribute INIT_31 of inst : label is "905D277B7760575247DCD261D3750C51524844911265D0B3489242741507384C";
    attribute INIT_32 of inst : label is "2209D0471582CDE4091849273491284426453709DDD27D249F4941B406868150";
    attribute INIT_33 of inst : label is "64D5CD5366745D09D17722511668CD0095A323404DD17102478911D24B5742CD";
    attribute INIT_34 of inst : label is "415534DE044C8245460915DCD103164520B32320C6235068060DD85AD26341C3";
    attribute INIT_35 of inst : label is "24D170A246645F645C051710991D955357436495052710D9C63014241778A247";
    attribute INIT_36 of inst : label is "742019D5C20911772241C6443445D8F4E467984C317D13745CD3645E28919381";
    attribute INIT_37 of inst : label is "95C944D16946440E34960B24587C19F3149C037254991D955355254669459245";
    attribute INIT_38 of inst : label is "665419D15D07166336474554DD0D58091031436684D0193D19C3045D366095D1";
    attribute INIT_39 of inst : label is "8937434096D9D1034593645746757151AD919DD5D98951DD99D500E55B152677";
    attribute INIT_3A of inst : label is "6CFDE79310748E689C61D47DFAA6F6736154D49C9D8C37D367D254F494D6820D";
    attribute INIT_3B of inst : label is "895A3FEFD9A566068C384CC153064C1D105D8757593840CD7F5DB0CDBF3F445E";
    attribute INIT_3C of inst : label is "CFFA894A25AE88C34DCA6A25370D2AB6BE166278E674D3F688D2630C30A6C86A";
    attribute INIT_3D of inst : label is "EA72530F3B9B2878C81AEFA384F32433BEF6177892197D2C38B22B0A8C3CB223";
    attribute INIT_3E of inst : label is "1126185551905102C3B7BF30E373734E3C3D30E30E8DBAB0F6EBDCEDD7CE4D37";
    attribute INIT_3F of inst : label is "0D04D134040554454D100D111D0CC345853340645CA904511013404434490410";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "E0268BA24DC2302909696664128248DA9A5432252C212FFFC22334488CCB0098";
    attribute INIT_01 of inst : label is "43234881303E40C0C4441CE860A4E0C3620C098410D902408C033012CE9204C1";
    attribute INIT_02 of inst : label is "E8300540B8B2002C9B2BB29240900BB8021124E8693844B0EC0A334234EE38D2";
    attribute INIT_03 of inst : label is "80792030CE028340F2030C3C8F08447D83123C344D213A0B4429B442A40C1C44";
    attribute INIT_04 of inst : label is "9202D98C0262C8009225A54E7E5A3009020A0038223B2030B4F93C05F00240B4";
    attribute INIT_05 of inst : label is "4F93C05E6409A2E6AA422480B665205920245599664B6992A05E90C112776744";
    attribute INIT_06 of inst : label is "404689A59440012955E118A212044AD5120020097E43CFA8F63CF900D3F4F027";
    attribute INIT_07 of inst : label is "125202A134F93C802A639F4208468C84048080C114460CA420296E9694C52221";
    attribute INIT_08 of inst : label is "94C00357DD23040B329D1030C492A5541059040948009544410511040816885E";
    attribute INIT_09 of inst : label is "A7B6A6273A665256125A6A562124102421784809080A10045A96A12C5154170A";
    attribute INIT_0A of inst : label is "00D0000000C000FFFF540F04FFF3AAAE55593004EF000228E840965699A62597";
    attribute INIT_0B of inst : label is "00F40100A047D08000F01400000540C000D0002A001FF4F800FD553FF0FF0080";
    attribute INIT_0C of inst : label is "F4F8F4FD57FFCFFFFFFC3F8FFDD2FC5FFFCABF3FCF3FC33FFF3FC300005050A0";
    attribute INIT_0D of inst : label is "551FD53003FFFF5053A3FFF4A9FDA367D387FFF296FFFF854BC757D2EA2A3F1F";
    attribute INIT_0E of inst : label is "005A5005A50055500154000000C04004055AAED26C65AA59048A4041412F3C15";
    attribute INIT_0F of inst : label is "F38FC2F0D62F9808BFFFFCFFF7800FFBFF6484C48EBF40A99800000015400555";
    attribute INIT_10 of inst : label is "54137FCAF813717CA723F06729C88C1CD5CA720FC07B28D815031C70410D07FF";
    attribute INIT_11 of inst : label is "FB8E3C8AA9300FC03C33645371080C0483FF0FC0385314C8605F1B1E36E49C20";
    attribute INIT_12 of inst : label is "443E1B4D130C3F94525AE8A172AE8A0A157C30CA05B744652FA60ACA87046182";
    attribute INIT_13 of inst : label is "2008B2702020080F1A3C5844103CA3E100C838C03E0E8003E0E8C2A3D20008E0";
    attribute INIT_14 of inst : label is "9180088A24B5480A428E323998AA66A98AAAA213A4C0A8E924B480D250C24600";
    attribute INIT_15 of inst : label is "4D234821418172208A59A4962789E26892782227F9375288F829E06420221430";
    attribute INIT_16 of inst : label is "830E838AE8AC2E3C3CA4A8F8A8FEA332021880525AD8883FEB858880E14E1C00";
    attribute INIT_17 of inst : label is "42892344C102344E8D005430C9C08620332348E20204130D2D222943BA2B0B8F";
    attribute INIT_18 of inst : label is "492402032D56594A509694999816B0032275674AD44225F59A6A293266006032";
    attribute INIT_19 of inst : label is "48C2C30F23C8090A3CA4AA4A906E30202523003280488429B4232030F802F24D";
    attribute INIT_1A of inst : label is "AE459030C32CFD3E520CF41F89138955D00912C1101540848184055FC64B0C06";
    attribute INIT_1B of inst : label is "4A44814DDC90D1603AC8D290831C30F069398B3030D2C2C342C3C3CF43CFC228";
    attribute INIT_1C of inst : label is "2A17FC3FE1344141E23408441D0246D8DE20B746073A1F869457DD680509B17F";
    attribute INIT_1D of inst : label is "80157CD61585CE07D530B4A2D4B65AD53B064A9A60267F67391B6986CEA8054A";
    attribute INIT_1E of inst : label is "1293BE92125C9E29A41CE10851FA681B9F9629E128E145F427F4174D2DDDAA34";
    attribute INIT_1F of inst : label is "DCF38734E181024D02D4E1C64D46D0A1D61C126090762842391F86B6457DDED2";
    attribute INIT_20 of inst : label is "66D0759401D4E7E1A12515F75A0111826C5FD101544D618EC7D537B4830B7346";
    attribute INIT_21 of inst : label is "0DC213C0618B02D194846B744847E18A815028D1F74488086491B50416662B90";
    attribute INIT_22 of inst : label is "9E110641B070AED3C4870451860A18B061863C1860B50180B708F1218646D06D";
    attribute INIT_23 of inst : label is "28DA278685E1B34AED4D67A909E1F278701CD418079010D4D67D71B59F951A46";
    attribute INIT_24 of inst : label is "2C191C4061CA3689E1A17860D8D40D67AEC1D359EC6DA6178709E1F04AED4187";
    attribute INIT_25 of inst : label is "068B1DC1DC193D06906734BDAA2D202C2EDA46A45D65445047EE518629D88B55";
    attribute INIT_26 of inst : label is "82A54518104074101D2C777637770C1DDD8DDD8BB0C10148474B74A4E617E43E";
    attribute INIT_27 of inst : label is "44076147520A10899CC1B250AED00C8860845060495297A8BAAA0B9714522AAA";
    attribute INIT_28 of inst : label is "95354D5254E2B91561946698AE45185507025491626956954165545D85CD95A9";
    attribute INIT_29 of inst : label is "D4D8414C75CE4107C099FD6C1D911D226660404410118812844B844BA1055254";
    attribute INIT_2A of inst : label is "87B1A5CED2D410160374B50535C2412904AC141732A2866069634B6040636AA1";
    attribute INIT_2B of inst : label is "937ACD41C2D6005062B5C2412904AC141C6D739074B5045CE412904AC14D7220";
    attribute INIT_2C of inst : label is "F6424ED9FA00B70808A019CA942614C0E6C1AAA11211D1DAAD7390760B5CE4D2";
    attribute INIT_2D of inst : label is "90B41B3A7183BA6807535F206986061F64686988293A390B51A2B083A2B50729";
    attribute INIT_2E of inst : label is "364AA4A0DDD4AA4A0D376D41376DC1C2DDA4267E2806A8E4EE80763A742A2A62";
    attribute INIT_2F of inst : label is "060267C55FD121D281D7C85FD8A98D14A4AE9899ADA6AAD82437AD8AE4DAD2B9";
    attribute INIT_30 of inst : label is "D2D7C95FB6AD804150A6D8E66AD805F67F4B7392B494E9253A616681942D5523";
    attribute INIT_31 of inst : label is "64267C647850B427D46517ED8A6363D2D7E485F217E29A526A63B0A69DF40763";
    attribute INIT_32 of inst : label is "A9829A75377D019ADF5B6AD805F2D0DAE66AD81F1A1253A494E9859A154D02D0";
    attribute INIT_33 of inst : label is "368DD81A0762D81188637060046488A1119372025E5596B7C55F21E7E54A6949";
    attribute INIT_34 of inst : label is "8212B8290005BC484AF12158836B367930A3256F0C22341091885C1A67EA223A";
    attribute INIT_35 of inst : label is "382096414967D28AD5C10910E12E112B86038421C10910E15D9025262564BC4B";
    attribute INIT_36 of inst : label is "660055D55E03D0E520C30D407B569818CCAB3805934AD4A5A5D4B5A590525142";
    attribute INIT_37 of inst : label is "D20B45F5E0474B4EC5FDF41498A0253C0424C3944A112E112B84144869499175";
    attribute INIT_38 of inst : label is "84462DE111880452344B844AE1C1144D1CC270A640E4193329C0357D6F7092D2";
    attribute INIT_39 of inst : label is "86984391F45992FF57D6D55747444FD29D12DED1E10D12DED1E1887C64252A77";
    attribute INIT_3A of inst : label is "D6DEDDBFB6FEE74F75FB9EBDF0DBACF2418AE49CE5009529652A7F4A981D0D41";
    attribute INIT_3B of inst : label is "4DFDB7CFF30F0D8C4C30E8C3030E0C3035F74F6E33BCE0CC373C7CFE3BBB6D3D";
    attribute INIT_3C of inst : label is "CDF3EE2F31C6E0D3CFD33FB8BBAE3BD0FF33836D74BCF3B8C4C3930C30C7DF2C";
    attribute INIT_3D of inst : label is "33E3930C3BCF783CDC0C72E0C0F378B0CCC7C3F5DBED6C3030F7C3CCCC38EFBB";
    attribute INIT_3E of inst : label is "28204455E52C290DC3FE3430E3C393CC3C3B30C30F0CB936CCC35F6CD30E4F3F";
    attribute INIT_3F of inst : label is "2DA0E4B4B497552DCE48A1212824538D903304D8DCDD1ED240038349304B12D8";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "2B45495A265AA9461465191B4052574E65188B45AC8B475DEA8BC2266D180CAB";
    attribute INIT_01 of inst : label is "F887ADF0AA3B0AAB2A7023074B090B05ABAA1E2E024C2B0AA9A4984A30EB4260";
    attribute INIT_02 of inst : label is "0F8A60E90D342242952150CB0AC331532A94A7034E348AB62D808AABFAB37242";
    attribute INIT_03 of inst : label is "0E34B545A61258E63B58698EE8048A84D8B434321428A849A2E42A226AA6B2A3";
    attribute INIT_04 of inst : label is "8232AA66B634D3AE86A2401C6E24B8D398D0B9D0B9D38A98A0E83A6215240A3D";
    attribute INIT_05 of inst : label is "0E83A6200028AAE28AA8A08CAA9825A82323A882A20A9A82AB8EAA698EA2A2A2";
    attribute INIT_06 of inst : label is "86292CEA72A22B8A8A68A4B4B8AAE0A882AE9AE86CA30EF8C238C88A83A0E98A";
    attribute INIT_07 of inst : label is "82B96AA9A0E83A69821F1B68AAE629222D242EEA62E6290D2908ACA02AE82AAA";
    attribute INIT_08 of inst : label is "5D4AA810A2BBE2658C6AABBE26640AADA9A36A4A08A72A22DA9A8B6A49A3AA86";
    attribute INIT_09 of inst : label is "9191925A519985995D0919122B4DA926AA1A2AD34A40ECAEACA076CEBA204DF5";
    attribute INIT_0A of inst : label is "004000C0000000FFFF55FA55AA04AA00AA009A005500B505C5724A4E44699291";
    attribute INIT_0B of inst : label is "0250008BE00050F02840000A800000F83840003F800000FEAAF400FF003FF0E0";
    attribute INIT_0C of inst : label is "ABFEABF4F8FC3FFFFFFFCFE1FC4FFEC57FAFFF304300FF00C330FFA0A00000F8";
    attribute INIT_0D of inst : label is "AA01F83FFFA0A3FFFFF85653FF9BE3FE53F1694BFF4A87FFFFF8384FFF3F87EA";
    attribute INIT_0E of inst : label is "00000000000000000000000000C900900FF00B14ECCF0000001000000030032A";
    attribute INIT_0F of inst : label is "002A08020104FFA8955401154001554101042A024410EF550900000000000000";
    attribute INIT_10 of inst : label is "0500C00E0A404840E62402503BBA4182040E62900944398A546480045161B155";
    attribute INIT_11 of inst : label is "1BECB24AAAFA5A003C3250100141411150882223821004000010801000024092";
    attribute INIT_12 of inst : label is "320AC3AAA9A2A061406B269982B266AC51A2BA2AA0A22233436765EEA8AA9A60";
    attribute INIT_13 of inst : label is "A9A68A8349A9A6908E4A0AA94A419484A40121290E491690249162ACAABA6B26";
    attribute INIT_14 of inst : label is "0D0A6AAA90910AFCDC308AC467B919043B42A99C26D80F0990AAAA4242903429";
    attribute INIT_15 of inst : label is "E9AEEF0A1EE982BA5075965527411244118C8B467BB842D1D6242FCDC9AB90A4";
    attribute INIT_16 of inst : label is "000800092BC9CE3E340D2CF104DAA489A8A2AA406B22A298A32A2AABCA5CEBAA";
    attribute INIT_17 of inst : label is "2CD0E129CAA8BA10FEA6068A2A2AA8A9ACBA639B5EA2AA20602B804248C0438F";
    attribute INIT_18 of inst : label is "2888AEDEA00920108C0B250278D8A5DEA8080AE90A69A19286282A8A2123428A";
    attribute INIT_19 of inst : label is "0AA90B8C232870C0339D2E106E829B76069AE802AE1AE302C96B94B8C636AA22";
    attribute INIT_1A of inst : label is "9C36A9079069C270B445F6B2EC8E60E06506B4D8CC802D2A2833200B030A6B83";
    attribute INIT_1B of inst : label is "AF21DB204904F41D3AE702CA5049048EB2789AEAEE029412D412D41E141E3024";
    attribute INIT_1C of inst : label is "404A08A0B8CAD436B849C1A1427030212B9C081151F0DB98492B20245852749C";
    attribute INIT_1D of inst : label is "A688AE0244343C76C1A681D206481526AC1C302C85026C8160D0B2B09C2458A0";
    attribute INIT_1E of inst : label is "460ACE0242212BA2C943B8C195B892439B8920E423B811B526E85AA022025050";
    attribute INIT_1F of inst : label is "2B2C1ACD063610127029067012B02106024948B1550AC194F0DB984892B20E02";
    attribute INIT_20 of inst : label is "8BFD80929421C6E614224AC8091644149D272A688BE0243C36C1A3A0AD40AC90";
    attribute INIT_21 of inst : label is "F29A6D05BC383024409912A901B8E680946F0B2D22920049A0840B51DA292705";
    attribute INIT_22 of inst : label is "0E4B5034F90C9CAD1218D1941942C38D0610D341840AC43C0843440650B02502";
    attribute INIT_23 of inst : label is "2900C39310E4F809CAB026E0F0E4F4393243AD48D1224BA5026C9C009B204C13";
    attribute INIT_24 of inst : label is "2242F1A5044A4030E4C4393207AB9026EE14FC09B70280C39350E4F909CAD491";
    attribute INIT_25 of inst : label is "513462E4A142C3512D08C950005F63E35E2412412022212236EE04D1020D1500";
    attribute INIT_26 of inst : label is "F5C0F265698D0A6142E10809C009FA420210024B2FA6162910080099E246CAC2";
    attribute INIT_27 of inst : label is "A0609D181FCBCBE00334F82C9CAEB2D248B30787A5A790A15003D781C9145400";
    attribute INIT_28 of inst : label is "AE9BA6EABAE2705A9AEA29A49C16AE2B2D8DA08EA402826A0608A1827850282E";
    attribute INIT_29 of inst : label is "2C3E36C10BEE3676E409B0264084402A292A0E2AA18A36826A0B2A0B1A56EABA";
    attribute INIT_2A of inst : label is "1B851BEE0423656F8C800850CBE21424D0B3476FB4B29B2546F8008D95842244";
    attribute INIT_2B of inst : label is "4C393076B22F850D8C8BE2142CD093476B22FB8D820851BEE142CD093472FB43";
    attribute INIT_2C of inst : label is "C218382FCE8E88E1E3B162B06D026D218F062EC44246060002FB8508C8BEE102";
    attribute INIT_2D of inst : label is "8D8878D1849C0B2C5894BCEF0630D0BCE183825951D0486294AD1CBD0529DBD3";
    attribute INIT_2E of inst : label is "CBD2C102A00D2C102A9096F690B6363220A1026EE458B58386C58AC1807BC184";
    attribute INIT_2F of inst : label is "10F026591B2406063606491B032032A0A09CA1A8024BF2B8E8809249C32D0270";
    attribute INIT_30 of inst : label is "0026491B892B8DA5AC8B2C229E88D1906C209D0D0A89FAA27685A27659D26CB0";
    attribute INIT_31 of inst : label is "03026589398D81F651B646E0300CB0002648199246E2240490A70C0B08A0D8B0";
    attribute INIT_32 of inst : label is "42302C094A28362C196892B8D992212C229E88594E6A27EA89DA3689DB229A2B";
    attribute INIT_33 of inst : label is "48122160580C0364310CADA7D1B2330446C80CC81304DB06589924E6C8089012";
    attribute INIT_34 of inst : label is "0F8270BCA106D20A0B482861D8015B8EA2E8D1B41B9CCA612611214026E0CBC0";
    attribute INIT_35 of inst : label is "2C92D98D01B8074926382C54982CA8272B22689AB82C749A66CA685051B2D20B";
    attribute INIT_36 of inst : label is "0842CE4E6B90240B445372904491216E6001A106C81F06C17606C1744140698D";
    attribute INIT_37 of inst : label is "02D265144B310BAB11BAA8DA88B606E0E0B1125A09A82CA827295A0A0AF46B0B";
    attribute INIT_38 of inst : label is "AA29A8EE8A68E284620B3A09CA38A158EC0D0419A1C3EE98C6E8598250A24206";
    attribute INIT_39 of inst : label is "10893F3DB60842D01A05B3B1B2A29C0248828CA8CA78828CA8CA97B79BD2C1A3";
    attribute INIT_3A of inst : label is "C1CCCD7CF9E0E39D3CD38E3C34E38D090409C1A3821A8274A27EB49DA3681836";
    attribute INIT_3B of inst : label is "0D3D334DD3CE0E0E4D30D4C3530C4C3135C31F1D3C30E0CC373534DD37733D30";
    attribute INIT_3C of inst : label is "4CD3DF0C30F0E4D30CD38D74770D30C0C303D34E3D34D334E4C3434C30DB2C0C";
    attribute INIT_3D of inst : label is "03D3C34D330E3930CE4F39D4D0C33135C0D3C330F30F1C3834D7534D0C34C703";
    attribute INIT_3E of inst : label is "08427B64E4210624C3343534D303030C3D3C30C34E0F783CE0C7CD0CC34C0C33";
    attribute INIT_3F of inst : label is "9203C702D25091C03C72A82C6CB2CB601CA7ED03230048007287691B7E30D46D";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "27298866200593F72611999B8F62666561988B369897F38EEA83D2220F6BF1BB";
    attribute INIT_01 of inst : label is "FB0FC883810B8A0A60E323333E7E39401B243E6C222E278A0825A08F33E7CE82";
    attribute INIT_02 of inst : label is "3FB202262FBFAA89662464E789E03C633648F3333E08C97C2F218207FC87CD2A";
    attribute INIT_03 of inst : label is "CE08BE38923862E8BBE38A266108CAD2FB330822F2AB08C0AC106AC52A4E9603";
    attribute INIT_04 of inst : label is "AA309A247EFEFCA8A261223F1A1278CF98ECA8CCB8EF8990A82A0A022200062C";
    attribute INIT_05 of inst : label is "82A0A020001A4BA0429A2A8C268A23AAA320AA82AA424AA003A8A64A0EAAAAA8";
    attribute INIT_06 of inst : label is "CAA45E5A3A92290AA92A90BF90AA40AAA264B2CA1890830820083909A0A8280A";
    attribute INIT_07 of inst : label is "A2A3DF9A282A0AC81A8FC62816425FEC2CAA6A07EE422CBE2A998BA82A0A2592";
    attribute INIT_08 of inst : label is "508AABFF869BC220E42829BC223DFABE2AAF8AAA98BDEAECE2AAB38AA8A9A4A2";
    attribute INIT_09 of inst : label is "98989BDBCD9DCDDD99A9899A272E2AA2928A99FF8A90E8A4B0A9BEBEA2A88005";
    attribute INIT_0A of inst : label is "AA0000EFE00000FFFF000000000000000000000000007FF6D6626A6266E81A99";
    attribute INIT_0B of inst : label is "FF0000FFE80000FEFF0000BDB80000FFFF0000FF780000FFFF0000FFF00000FE";
    attribute INIT_0C of inst : label is "FFFFFFABFEFFCFFFFFAAAFFEAAFFFFEFE7FFFF1555155515550414FEFA0000FF";
    attribute INIT_0D of inst : label is "FF15550554FEFAFFFFFFFFFFFFFFE9FFFFFEFFFFFFBDB8FFFFFFFFFFFFFF78FF";
    attribute INIT_0E of inst : label is "00000000000000000000000000E002000FF00F00FCCF0000000000000005543F";
    attribute INIT_0F of inst : label is "0FEAFBFEFFF0AAAB800001403FFFF01414FFEAFEF14020550800000000000000";
    attribute INIT_10 of inst : label is "FFFC000AFAFFFBFCAEEFFEFF2AAAFFBEFFCAEEBFFBFC2BBAFFEFBFC0FFEFAC00";
    attribute INIT_11 of inst : label is "8BCE38D664FC81003C308055554555155111044014551545545515553FFEFFBE";
    attribute INIT_12 of inst : label is "3329EFC82AA06D33292864A2A28646C4CCAC92C9088888BBEBAE26E68B38D302";
    attribute INIT_13 of inst : label is "29A0B2537828A0620C88808CED88488ED8A623B620843362884332A5829A0968";
    attribute INIT_14 of inst : label is "CDEA0A2A088889E3E333825210C484020C9A680CE4F21F3908A0A6222AF73728";
    attribute INIT_15 of inst : label is "A90A433232B2A2B1FF28A28A22A0A23A0A888B31B9AD22CCE2220E3E382888BD";
    attribute INIT_16 of inst : label is "C614060402323409093F30323822A18193A8AA292868AE46574A8AA3F23F2824";
    attribute INIT_17 of inst : label is "8EFCEF2FF8182C33FF2022B20A64AA2AA1B242B30A42A2CA2A247C85009C9D02";
    attribute INIT_18 of inst : label is "2908840084843330CCCC23213800940080888A8B4A8B28628A950A82A2A37282";
    attribute INIT_19 of inst : label is "8A4A48822088CC9E084F332322A6ABAC92A24462AA3AA33308EA8C8826308A42";
    attribute INIT_1A of inst : label is "4D0064208208E238B308E2B6CB0AC2A2A2327FF0C8889FEA8A32222A4B8A090B";
    attribute INIT_1B of inst : label is "92C2B2CAAF30BCCC2FE3A2B102082081C22802A0ACA230C230C230CE70CE6B90";
    attribute INIT_1C of inst : label is "AE8A5A2590C9B31090C88C9F33E33323290CC88404FCC68608A2221000CE2288";
    attribute INIT_1D of inst : label is "B9C8EC2021013F3188A0A822A1AA86A2653F3330A3301888FCCCC2272310009E";
    attribute INIT_1E of inst : label is "22261E22222029232F3290CC8C6848CD068422E2269088674198099A1AA92E88";
    attribute INIT_1F of inst : label is "2A68CA9A3202F3C0F32232F300F32632201C14823CCF8C8CFCC6860C8A222E22";
    attribute INIT_20 of inst : label is "18840809F333F1A1822228888400333388A2279C8E02023F31889998AECCA9B3";
    attribute INIT_21 of inst : label is "F2F029443CE52323820869D880A982A2812B3B2B5D8810C0988CC805C9941340";
    attribute INIT_22 of inst : label is "2427CE01988E4D69480A04A8CACECE5A3233968C8CCBFCCCC8CE5282F3F32332";
    attribute INIT_23 of inst : label is "2F38CD06334398A4D62301A233418CD0E2276F3FC722276230188CC806223886";
    attribute INIT_24 of inst : label is "222294ACF18BCF33418CD0E223622301A40188C0633289CD06734398A4D6B3C6";
    attribute INIT_25 of inst : label is "C7AD33E26332A7C7CCC8C820000BF3C30A1231202203233201A42386822FC222";
    attribute INIT_26 of inst : label is "F0B332332488C9223284888B8C84E422222321074E43022888888A48A02189A7";
    attribute INIT_27 of inst : label is "989C80488C2C82422741989E4D6920CD889DCDCDD0A2881C2557C2CCC8CE0955";
    attribute INIT_28 of inst : label is "6A0A82A1A8C13401471994504D00711AC90C988DACE2611989E6627236332631";
    attribute INIT_29 of inst : label is "286832848A8E32018CC06222226222259425C99572650169198759874602A1A8";
    attribute INIT_2A of inst : label is "8B88CA8E2027272A0C8A088CCA823310CCC3332A3E028C2232A0909C9CBCE122";
    attribute INIT_2B of inst : label is "0CF43332302A08CC8C0A823330CC43332302A38C88088CA8E3330CC43332A3C3";
    attribute INIT_2C of inst : label is "127F3F321E4C08CCCCC0022327302B53FA4CE3222222222552A388C8C0A8E331";
    attribute INIT_2D of inst : label is "8C09FB8C9C9CCC700080A1EE32332361E23231389C9CF89D8C88CC88C8D8088E";
    attribute INIT_2E of inst : label is "0CF33232622F3323264842C248C2023022E3301A1000C3333300088C88FA8C8C";
    attribute INIT_2F of inst : label is "3333018886224222102188862AE2AA58984D60660108C26C18884104D0322134";
    attribute INIT_30 of inst : label is "24218886842380ACAC0C28594E080860188088C9C968C65A1180A03088222929";
    attribute INIT_31 of inst : label is "37301888A08C0821882221A2ACAAA1282189086221A110CC40CFCCCC261808A1";
    attribute INIT_32 of inst : label is "0333308A098602284628423808622D08594E08062C25A31968460280CA433027";
    attribute INIT_33 of inst : label is "8BA22A2A88AB2A22ACA88CBB8CA03AF222809E8886218A118886228188844331";
    attribute INIT_34 of inst : label is "426134281332A5A98A962622B2A8CA1A2CB18CAD2B0EA933333B232001AAB69E";
    attribute INIT_35 of inst : label is "082088C0A4A1A084A2A708E8361D66135A4098262708C83623B2D8CC8CA8A587";
    attribute INIT_36 of inst : label is "88CDAAAA2B02208BF0823A33188623093904E332B282A1A862A1A863302924C2";
    attribute INIT_37 of inst : label is "A2FC886189988AC94866180960AC92A49C2320C9A4661D66135809898623268A";
    attribute INIT_38 of inst : label is "5894E2D221399C8D8D874984D26323632B48D8C8D3F3280E4290C86A1AAC22A2";
    attribute INIT_39 of inst : label is "33808FCC6226228686A1AAAA888882A232222D22D232222D22D22A8D88CECC8B";
    attribute INIT_3A of inst : label is "A0CCCA24689082082CB2890920A2090488C4D06232E7CA109A31A18460263602";
    attribute INIT_3B of inst : label is "082C330CC2CB0B0B0C30B0C2C30B0C2C2CB2CA0B2830A0CC332830CC33330A28";
    attribute INIT_3C of inst : label is "0CC2490A289090C30CC24924330C2490924202892030C33080C2030C30820808";
    attribute INIT_3D of inst : label is "02C2C30C330B2C30CB0B2CB0B0C32C24B0928220B2CA0C2830A2830A0C30A283";
    attribute INIT_3E of inst : label is "3C92A32AAA633229C3242430C242430C202030C3080820208092080CC3080C32";
    attribute INIT_3F of inst : label is "42F3FAC90928AAB23FAD5222692CB2CA28BECE1322128B28A24AC49BAC3CEFAF";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
