-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.Vcomponents.all;

entity COSMIC_ROM is
  port (
    CLK  : in  std_logic;
    ENA  : in  std_logic;
    ADDR : in  std_logic_vector(12 downto 0);
    DATA : out std_logic_vector(7 downto 0)
    );
end;

architecture RTL of COSMIC_ROM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'    => result(i*4+3 downto i*4) := x"0";
        when '1'    => result(i*4+3 downto i*4) := x"1";
        when '2'    => result(i*4+3 downto i*4) := x"2";
        when '3'    => result(i*4+3 downto i*4) := x"3";
        when '4'    => result(i*4+3 downto i*4) := x"4";
        when '5'    => result(i*4+3 downto i*4) := x"5";
        when '6'    => result(i*4+3 downto i*4) := x"6";
        when '7'    => result(i*4+3 downto i*4) := x"7";
        when '8'    => result(i*4+3 downto i*4) := x"8";
        when '9'    => result(i*4+3 downto i*4) := x"9";
        when 'A'    => result(i*4+3 downto i*4) := x"A";
        when 'B'    => result(i*4+3 downto i*4) := x"B";
        when 'C'    => result(i*4+3 downto i*4) := x"C";
        when 'D'    => result(i*4+3 downto i*4) := x"D";
        when 'E'    => result(i*4+3 downto i*4) := x"E";
        when 'F'    => result(i*4+3 downto i*4) := x"F";
        when others => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO   : out std_logic_vector (1 downto 0);
      ADDR : in  std_logic_vector (12 downto 0);
      CLK  : in  std_logic;
      DI   : in  std_logic_vector (1 downto 0);
      EN   : in  std_logic;
      SSR  : in  std_logic;
      WE   : in  std_logic
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
    rom_addr              <= (others => '0');
    rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "554464B24000841DD9594759C74C20D915508454610C6118600001294201B113";
    attribute INIT_01 of inst : label is "355C449DAA23347547745108046AAAAAAAAAA0192376892E80020415551D4105";
    attribute INIT_02 of inst : label is "220620021F61F61F61F6185D86176185D8617410086D0AAAD70008414D244378";
    attribute INIT_03 of inst : label is "D2410491413491654765474575744646445478B61B61B61B61D800888A28A28A";
    attribute INIT_04 of inst : label is "1D34C34012341351C641476165CCD56D05478808054765451524451144934924";
    attribute INIT_05 of inst : label is "244889AA0255B45620014417191E746A1B8956446013055B8E134104D3544D47";
    attribute INIT_06 of inst : label is "06788110519D9D04465547013404D344D471D0C042D041104015075A84807341";
    attribute INIT_07 of inst : label is "8681E059055544000009B15FFE943E9051510C102035CD048CC803215B35590E";
    attribute INIT_08 of inst : label is "706520756074411025CFFAF50F5308510461441103206A9433046681E4690668";
    attribute INIT_09 of inst : label is "1209C06120A2242224104248424AC270016450C1468000D07309C04355249530";
    attribute INIT_0A of inst : label is "424515066256140514991411C34826045C1449C3482625564535734462449C00";
    attribute INIT_0B of inst : label is "5002382A404D501500E20801501591576642046341E0A0014040270000000000";
    attribute INIT_0C of inst : label is "AAA07455011A050459056050601826416082C240207302281502A206049C134A";
    attribute INIT_0D of inst : label is "670654981074CD04009E0C074276140414524A16B4DC26A241B059076CA41905";
    attribute INIT_0E of inst : label is "D042C278800DD3400214D047344B270800D14D4342011C3B0D026CC0023441D1";
    attribute INIT_0F of inst : label is "80572360DC858153749C0216044908091374210DC240004507706420D343811C";
    attribute INIT_10 of inst : label is "144466554465544742254201460007413310E4DF804504518D130D1D11410420";
    attribute INIT_11 of inst : label is "0190904CC01E90890D4D107A4324352A86344274912686817174C511595511D3";
    attribute INIT_12 of inst : label is "480D542000551545515481D5B3365003450567454D147057448220E91D208800";
    attribute INIT_13 of inst : label is "D0CE04744C4448012511DC004D141645520AC01B6582B7419EBAE84CD162511D";
    attribute INIT_14 of inst : label is "6412034525388412035D00030066666620C005145140448017494E080B81305C";
    attribute INIT_15 of inst : label is "52001442098250526488381585010198585C15E074C44480D98D52480D760563";
    attribute INIT_16 of inst : label is "0CE000000000000000000000285591D1185591D180051059C4771052D50D15A1";
    attribute INIT_17 of inst : label is "5420014714447710A753700017D1451144147477905504CCC2394D924A179E20";
    attribute INIT_18 of inst : label is "2BA8EE536492B88800510182200144060C30398805116DC20014714474418948";
    attribute INIT_19 of inst : label is "000F5D64EC00DE84880D5810110081100221A064123241054201064101054082";
    attribute INIT_1A of inst : label is "727245B28611504705525430D1D10413895264D18611C21223110E00FA50F900";
    attribute INIT_1B of inst : label is "56E05DEE80016110E591AB45B01536DCC005914D94D3405D128D1D1115114930";
    attribute INIT_1C of inst : label is "4E0916C156B44A347444544531448518591AB6CC0A00156CA510D5802D5B45CB";
    attribute INIT_1D of inst : label is "000000053852C53B83E7C2513C033029127855241B46CE1AB64144499051C1B5";
    attribute INIT_1E of inst : label is "95D3705D3609D1192781192405246141745185099D5910D191E34991480D8354";
    attribute INIT_1F of inst : label is "00C062012422012416012437C5D994DDCD96134D02402660917605341CE851DD";
    attribute INIT_20 of inst : label is "5768585A28601941019107764D9526983763640DA645DC59494535A49515850D";
    attribute INIT_21 of inst : label is "1F41F71F61B51441042A9555554000001B222222222222051344434A946A9051";
    attribute INIT_22 of inst : label is "544105554748A55464A01D7654044B9AE04516B84A594641555167A74C21F601";
    attribute INIT_23 of inst : label is "400AAA9FFFFC03FFFF9554553655587FE00521E007F1640415551D5501055547";
    attribute INIT_24 of inst : label is "C7C711100A4A410113807FC438110AA400AA4113FC4007FC1100040040012AAA";
    attribute INIT_25 of inst : label is "7F310041F1C40110041010401100410104011004AA904012AAA7F2AAA91C7C40";
    attribute INIT_26 of inst : label is "110AA410AA41107C4107C411040AAA404110407FC40412AAA900AAA91FC72AA4";
    attribute INIT_27 of inst : label is "89924D93491024928534145222088E4E2AAAAAAAAA91FFC71C7FF11000410400";
    attribute INIT_28 of inst : label is "4524345309D24455D47194924A3351C445247091490514C2749114751C552410";
    attribute INIT_29 of inst : label is "C9930D04DD0634D80701245092645D8926455892601E43000448230D1D471DC2";
    attribute INIT_2A of inst : label is "7193093442080DC50E60D20D55349146145424C00080000D1002B4D050D34411";
    attribute INIT_2B of inst : label is "10B8CC0FC0CCB81000CD471D80D500C0157045046176AA81120D5244510491D7";
    attribute INIT_2C of inst : label is "AA80B24404081D767657656C81576571771C80536371171C6401341B73836400";
    attribute INIT_2D of inst : label is "3FC02BFFC03FFF4000002BFFC000003FF82AAAAAAAAAAAA9B35F214C933060D2";
    attribute INIT_2E of inst : label is "C01FFFC0003E80003FC00002FFFE80003FF8003FC00002C03FC0383FC002C000";
    attribute INIT_2F of inst : label is "000000003FC0003FC0080A8CFC2A0203F3002BFFC03E80003FC02BC03FFE803F";
    attribute INIT_30 of inst : label is "450000014A00000A14000000504000105000000014000001400000000A00000A";
    attribute INIT_31 of inst : label is "C00A00003E400A1FC00000003E40001FC03C00D4507003D0514A008514200A01";
    attribute INIT_32 of inst : label is "FC0018003FCC083FCA80000FFC00000008000A8D5F6A001F0F000A003E40001F";
    attribute INIT_33 of inst : label is "FF000002AC40003C5300AA8CCCE82014930000915FC0003D51000001BFC0A83F";
    attribute INIT_34 of inst : label is "004000400000000000400040000008000800003FC0000000FF00003FC0000000";
    attribute INIT_35 of inst : label is "0000001007C0001C9040000007C0001C90100050001000100050005000100000";
    attribute INIT_36 of inst : label is "400AAA1AAA5AAA5AAA5AAA7FFFFFFFE8002AAA802ABFFFC088101F5C90100000";
    attribute INIT_37 of inst : label is "57F557FFE7FFC3FFFFC000256000000000256025602560256005400540054005";
    attribute INIT_38 of inst : label is "02BFFFFFFFFFFFF555FF55FD75FFFD7D7DFD5F7F7FFD75F7F5F7FFFD55FFD5F5";
    attribute INIT_39 of inst : label is "0028002AAA802ABFFFC00020003FFFC000BFFFEAAABFFFEAAABE0002A83C0000";
    attribute INIT_3A of inst : label is "75D11621DB4518D584C55DDDE8D5912524410460445D146451074109160C5814";
    attribute INIT_3B of inst : label is "C915465938C91546593814C915465938274DD2549127206CED02010C5C02041D";
    attribute INIT_3C of inst : label is "3A404040CB10001A47A0F2432393913B93B555FFFFC420000000E64F91393938";
    attribute INIT_3D of inst : label is "E1C130A808040C92C133A804040C910041C2F4441C274B441CAE2211A324C309";
    attribute INIT_3E of inst : label is "0332B32B40379FB49068B0C344D10402F0500E20310B03303CD10402D1244B80";
    attribute INIT_3F of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAF1D9D9F99153B993999999333333";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C30C94614A028A2D6DA0C87A1F8870FE1F982FB8C120C318B00003364AAB0023";
    attribute INIT_01 of inst : label is "8761FA92AA3F14766564322AA1EAAAAAAAAAA3F6AEDA4AA987130A030C3E0280";
    attribute INIT_02 of inst : label is "3002F22A64AE6AE4A66A64A3B9AAEE6A3992AC1024AA0AAA0A6024A1C71CB14C";
    attribute INIT_03 of inst : label is "31CF1C33CF2CB2C4477776494476944774B48CBEB9E3BEB9E3E04892AD36D36D";
    attribute INIT_04 of inst : label is "7A8701E0F60828761EA1F48094C06112084A0B142D877747D23F83E0F870C33C";
    attribute INIT_05 of inst : label is "CCAC099902A6486A102080047612EA992440747662D21A660DD0823CB2E4A1C8";
    attribute INIT_06 of inst : label is "004882001E16120848585A0D083CB2CA1C87A802CB208B608966D82A88F01C82";
    attribute INIT_07 of inst : label is "4002DC8600000000000171C5555540001A1107B2001C7209C9C00A6044384722";
    attribute INIT_08 of inst : label is "8096019B619B47203CC005005511249248B2CB220127AABB8024A002DC864A00";
    attribute INIT_09 of inst : label is "25DA9C9B5C103B02090071D401C781C12388E0C0C344B0A04C0F8341C9187D30";
    attribute INIT_0A of inst : label is "B56DD5B56B96AB47D452DCD600F00F1B531F4380F00D1474761B71B471C87449";
    attribute INIT_0B of inst : label is "5120E4B943C35CF28D9C030DDBAD2387477F28B08A9EE437429027F000101002";
    attribute INIT_0C of inst : label is "AAA288E2CAAA8228E228A261C0A03C7A1FC703C42C5C1264E2EE602928E4A3AA";
    attribute INIT_0D of inst : label is "8B0B4AD862B8022800FA0828877809090AAB6A3A88A43EB08A6CE2289BD42D86";
    attribute INIT_0E of inst : label is "20C303E0448A22A13108A94B1955193848A24282BF8F2C0F0343DB0411288A23";
    attribute INIT_0F of inst : label is "83C93090A4064EDB4BA84A1B3B6DFC0F228A3D0303C122992B60B7F422834324";
    attribute INIT_10 of inst : label is "0784A56565565655701652116711154033018951B3C918F3C328252598A98F3E";
    attribute INIT_11 of inst : label is "00649AF00A096AB6C98E9825A8DB262AA6A484CB32A64300D09641E129999959";
    attribute INIT_12 of inst : label is "448AA8122829284A908429619C185023828845846E5985444448D25034D23400";
    attribute INIT_13 of inst : label is "241201440B044089015110080E08044471250897414145661596580B52501511";
    attribute INIT_14 of inst : label is "8411284609C448D122AE089B2291919100C08A082082444A184271C494802C70";
    attribute INIT_15 of inst : label is "C10208830F41E0B08484880202428A1CA0A0A12004BC400861C610848ABAFA91";
    attribute INIT_16 of inst : label is "850000000000000000000000241D1D12281D1D1240820016886A2A1A6D46D1A1";
    attribute INIT_17 of inst : label is "20CE208306886A2A8B4262222A2282208004A84AE8768F0143C44E13AA1EB108";
    attribute INIT_18 of inst : label is "2864111384EA8094082001925020800649C106808220AACCE208306868728244";
    attribute INIT_19 of inst : label is "0005500000E490E05003202420CEC20CFF0C405A112050286003086032286031";
    attribute INIT_1A of inst : label is "90A386CC470092B62B6294825259DE9A4761C83280925970131779FFAAAA5500";
    attribute INIT_1B of inst : label is "87B01E1108A093001161AB86CCF20F29448E238A2C2280F121E52592992A6DC2";
    attribute INIT_1C of inst : label is "A14E1B33C8448794964A64A980828204161ABB7801AA18731124E144B21CA18F";
    attribute INIT_1D of inst : label is "000000154104003FC17E640014082021684462BB0FC3B11ABBB19A86EC6282DC";
    attribute INIT_1E of inst : label is "29DB779DB607569DB7729DB7071C809074720241DDDDD8DAD2FF4BD2C802C280";
    attribute INIT_1F of inst : label is "A203860E861D0E861C0E861F01D1D06D46D1008A83C41C8071C8071FE5509955";
    attribute INIT_20 of inst : label is "CBA8B8BA2CB0A24242D02B756DD5B5550B60B40A5582DC2D42822856F5AF4E12";
    attribute INIT_21 of inst : label is "2AA2892A92A92092083FFFFFFFFFFFFFF7A78D278D278D01238460AA846A10B2";
    attribute INIT_22 of inst : label is "848280C30F8094F42E0A0F3D490A0F03C80C30F2494343E030C32C178CA2A902";
    attribute INIT_23 of inst : label is "80180062AAA400AAA94000014100001F009C40000EB0490A030C3A124280C30D";
    attribute INIT_24 of inst : label is "3EBEE614180181466001E4B80066181801818660AB8C1EA46600180180066001";
    attribute INIT_25 of inst : label is "EA060187AF58066018606180660186061806601860618066019EAE18067BEB80";
    attribute INIT_26 of inst : label is "66001861800661EB861EB86618186181866181EAB8186618180181867ABEE01F";
    attribute INIT_27 of inst : label is "C320C3E0CF280CF3C30E3C303E250FFA000000000007AABEFBEAAE6001861800";
    attribute INIT_28 of inst : label is "C33E2C32CF20C8321D8728A3CF2C761F8F3CA030CF8F0CB3C8320E8761DA3871";
    attribute INIT_29 of inst : label is "4229033CF29838F03D0F3C38F3D83E863C832823F0F50012C89702CB21C87AC0";
    attribute INIT_2A of inst : label is "8722C32CA1038B39719030C3220C33C908F80CB0EC040C0B244A88A05CB0C83E";
    attribute INIT_2B of inst : label is "FCA864098064A8FC00B1C87A885240D8F7B4492852B6AA46110320D8321CF21C";
    attribute INIT_2C of inst : label is "AA876D488C08966AD92E924C89E5AFBADBAC8966AEBEDB28409AA9A6B0C3F400";
    attribute INIT_2D of inst : label is "FF02FFCFF83FF4000002FFCFF800003FFFAAAAAAAAAAAAA937FC0A0104341212";
    attribute INIT_2E of inst : label is "C001FFC0003FF802FF00002FFFFFF802FF3F800FF8002FC2FF003F8FF82FC002";
    attribute INIT_2F of inst : label is "0000000027C0003D8001928630286400C902FFFFC03FF8003FC2FFC03FFFF83F";
    attribute INIT_30 of inst : label is "C003C0C005303C050000A080A0A0A020A00000003CC00033C000000005000005";
    attribute INIT_31 of inst : label is "5805800027C0253D8000A000A7C0A03DA000A080A0A0A020A00500403CD00533";
    attribute INIT_32 of inst : label is "F006042507C4903D2000B403FFC0002AFC02D147003D5800F9009500A7C02E3D";
    attribute INIT_33 of inst : label is "FD001F8117C20835F4092A8CC62186152401808001C0201000002B49FFDB833F";
    attribute INIT_34 of inst : label is "000000000000000000000000001EBC1EBC00381FE00B000BFD00381FE00B000B";
    attribute INIT_35 of inst : label is "00008080E7E0001D00008080E7E0001D00000000000000000000000000000000";
    attribute INIT_36 of inst : label is "A03000EAAA800A8A808A0A3FFFFFFFFC0007F54BFFDFFFC0FC022E5D000382A0";
    attribute INIT_37 of inst : label is "16F516FEAAFFCBFA8A800005400000256005400540054005402970263026603A";
    attribute INIT_38 of inst : label is "03FFFFFFFFFFFFF000F48A328A3FD2328E32A33000328A33CA315572A23A95F5";
    attribute INIT_39 of inst : label is "003C0007F54BFFDFFFC000300035554000D555D5557FFFD5FD3FE02FFFBC0000";
    attribute INIT_3A of inst : label is "3C32892AFCAD206DAA8A2D6DD8A2D2B628830CA3883E0C3C220F830F3A206884";
    attribute INIT_3B of inst : label is "C922CB3FC0C922CB3CD118C922CB3FE10A5324CB32A527BBC2022B3024880A0F";
    attribute INIT_3C of inst : label is "278B441CBE092705123CAB8042D45718043000FFFFE10100000242903D414140";
    attribute INIT_3D of inst : label is "F010437CB441CBC0104230B441CAD24C080A70FA80A7C63A028E3041C238441C";
    attribute INIT_3E of inst : label is "01CCDCCC00041CC0839F7CBF4B0041CCF084EF09043F40C3744041CEF151008C";
    attribute INIT_3F of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA72AAEF7A66E99A69AFA5FA9E94E9";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "1652B2EB2760462C2C21084A13B6A90243A601BEDB6041188C0003250AA80C89";
    attribute INIT_01 of inst : label is "44E11B02AA4090300001422AA6AAAAAAAAAAA90A442A12C2AC994B58698A7AD5";
    attribute INIT_02 of inst : label is "522934095DDDCD1CDDFD977F459ED557B455DCB6077F28008CB705671040BDAA";
    attribute INIT_03 of inst : label is "C71851441041043332222209110191100183AA51041C614510E900F3FDF65B5D";
    attribute INIT_04 of inst : label is "42ECF485A9AA244E12B4108C1B2D0EEA8B0A2AB640A11110424090E439C41061";
    attribute INIT_05 of inst : label is "6393120A943BAAE9B6024C82BE09F9EAB0080809FBAA53BA2AAAAE4104309128";
    attribute INIT_06 of inst : label is "87AE1C3206C0EA880B0B1A2AAA41040912842ED79CA89C6D0192667AB902B2A2";
    attribute INIT_07 of inst : label is "4230E473200000888884480000000002002B5C3622720A8AA0214087B2508A4B";
    attribute INIT_08 of inst : label is "14094C088C08902D6B200000000A44514491451A2B456AB489444230E4734423";
    attribute INIT_09 of inst : label is "9EE32667ECA4E2C0F0C1E4B6179C37B40140721492D014B2A0DA8AA40841298E";
    attribute INIT_0A of inst : label is "089202480BC0BD904140614274A241C1A8411214A241D8080B48B489E7290929";
    attribute INIT_0B of inst : label is "9404B97E1552B1521EE8902CE6BC01C0C0E754A413CAF0801985290595158515";
    attribute INIT_0C of inst : label is "AAA4485298AA504C524486D59535682B09D61680AAA0C3B952AF84C0C03500E3";
    attribute INIT_0D of inst : label is "48404B3504EA104C0055014488485850D2F4EA1E80B36AB413A05244A8338350";
    attribute INIT_0E of inst : label is "0492D6A2900902C330C0B809408AC2C900923032E7902550D656AC3022249121";
    attribute INIT_0F of inst : label is "56085C0CBB103C2CE8290040F0B39C9822486A5E76A4044850C60E7502CA9021";
    attribute INIT_10 of inst : label is "818190909080808084C094CC095CC08033023502440841A69CA890220BD2DA60";
    attribute INIT_11 of inst : label is "21A162C32816A68A3612705A9928D8401E90A6098E489655940AE0602424242B";
    attribute INIT_12 of inst : label is "D01D8CA4A09F07C5B06CAC22A0C8B700418831832F08CB0B0B2501502493EA1B";
    attribute INIT_13 of inst : label is "212B84A4DFB2B21E20E0EDC0410C838384AED0384F8B03960E38E0DFC2C20E0E";
    attribute INIT_14 of inst : label is "88B4A24329CB2834076329C24ABB57312294053C12CB2D2806CA72128AE17D21";
    attribute INIT_15 of inst : label is "BF602488DA94AE240AD2AE1212381C23854B02B86DFB2F21221222901D8E08C4";
    attribute INIT_16 of inst : label is "000E44E80000000028282828AA020202A6020202D809320EAC3A76E422122C04";
    attribute INIT_17 of inst : label is "02B3424D83883AF60AA6DE4027F34D224C80B81AF5021AD0F6880300E042F025";
    attribute INIT_18 of inst : label is "40AA2000C0380AAD4093208AB5034C82280C8A6D0D227F2B3424D83839025023";
    attribute INIT_19 of inst : label is "FA5000000000909000902323C3AE3C3AE7480C1B2CAC87E08417E08414C0852A";
    attribute INIT_1A of inst : label is "0D0C03AF128F070870BD0A890220BD2C902739CA0B0A0008C882320000000050";
    attribute INIT_1B of inst : label is "EE32CEECD0225D32E0600383AD0252F2900501C92302C98C249022022064BB0D";
    attribute INIT_1C of inst : label is "9E700EB40BB0924088088192EC8C923206003A056CAA07ABECA1CE9027C9DE38";
    attribute INIT_1D of inst : label is "AA0A0A800000003FC00000000028A5AC27B812EC19CE7E003AC04B34B01A909C";
    attribute INIT_1E of inst : label is "2C3FA0CECC56C2C3FA82CECC5650848439421210EC2C21C6CAA31EC7BA7072C2";
    attribute INIT_1F of inst : label is "7435C8D78959D7895AD7895A2030312312328C0B368A508D65085652BEE1CECC";
    attribute INIT_20 of inst : label is "0B01C9CA79C912143438D0C493124C0048C48DCB00523523B0B02C82F0BDC522";
    attribute INIT_21 of inst : label is "1DD1DD1DD1CD10D10C9555555555555567B8E38D34D249202FC09EE0080029C7";
    attribute INIT_22 of inst : label is "B0A2D61A62AD13F1FD2B545908496398ED61A63B913F1EF58698EC93A119DCF1";
    attribute INIT_23 of inst : label is "2A8000000002A80000BFFAFEAEFFF03901000008AFEB084B58698EC212D61A63";
    attribute INIT_24 of inst : label is "000000D7C0003D700D7C0003D700C003FC00300C0032C00300FFC3FC3FF00000";
    attribute INIT_25 of inst : label is "0000FC300003F00AC30F0C3A00AC30F0C3A00FC0000C3F00000000000000003F";
    attribute INIT_26 of inst : label is "00C0030C00300C0030C00300C3C0003C300C3C0003C3000000FC000000000000";
    attribute INIT_27 of inst : label is "900490C4902D4124904B41229515555500000000000000000000000FFC30C3FF";
    attribute INIT_28 of inst : label is "10494128102419061384E50492804E109040A50412504A04090E4184E1294124";
    attribute INIT_29 of inst : label is "1C25DE41024861274950412524290E1841902344A5250B4A66BB281021284214";
    attribute INIT_2A of inst : label is "84681040841010CF8CC524902049040B412549050E3C59D02D0280B2F107094E";
    attribute INIT_2B of inst : label is "A8A8A8CA8CA8A8A8FE012842184214C10DF80A408D3AAAD02290240906410213";
    attribute INIT_2C of inst : label is "AAA4E32F3CA91974677773229117447B777291D4447377322D15FDDFDAA438FC";
    attribute INIT_2D of inst : label is "F40FF401FFC0003FF80FF401FFFFFF40002AAAAAAAAAAAA84000BFE14586C856";
    attribute INIT_2E of inst : label is "C0000002FFC1FF3FF41FFFC00001FF3FF43FC001FFC03FFFF4003FC1FFFFC03F";
    attribute INIT_2F of inst : label is "00001BC0003E400000092FC2403F8600180FF43F4001FF001FCFF4003F41FF1F";
    attribute INIT_30 of inst : label is "0A000A03C0CA00303C0050405050501050003CC00033C00000000A00000A0000";
    attribute INIT_31 of inst : label is "89001BCA403E40001A005BC0503E5000500050405050501050003CCA00B3C020";
    attribute INIT_32 of inst : label is "40004BC0923E0A420603F0007FC0003FD0090001AF8A0621A401ABCB003E4502";
    attribute INIT_33 of inst : label is "D4022BC02F7AF80104024A8618463315490000C240C040006000F6CC1FFFF93D";
    attribute INIT_34 of inst : label is "000000000000000000000000000BFD4BFD403F07FFFF003FD4003F07FFFF003F";
    attribute INIT_35 of inst : label is "0000DBC0406E00100000DBC0406E001000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "40055500E92A90F430E050FFFFFFFFFC03C07E2FD407FFCF03C3415000011C4E";
    attribute INIT_37 of inst : label is "FFFD7DFE99F155354540002560000005402630266032603AA000501150101010";
    attribute INIT_38 of inst : label is "03DFFFDFFF7FFFF000F3CF33CF302F33CF33F33F34B3EF332F32A8B36F35F5F7";
    attribute INIT_39 of inst : label is "003C03C07E2FD407FFEAAABAAAB0002AAAC000C0003FFFCBD03FFE3FFFFC0000";
    attribute INIT_3A of inst : label is "59428B41DEEC214E89502C2EE102C67840904084090649214240924852B10FBE";
    attribute INIT_3B of inst : label is "9192673CCA9192673DC9C29192673CC9C09826098E4B457F22AA9703036C6B54";
    attribute INIT_3C of inst : label is "AF063A02AF3E908002B8E7495A1503E5503000FFFFC204000002954281555556";
    attribute INIT_3D of inst : label is "C3285A3C63A02BF3285AF863A02AD3C15150CC00150C844054320C080A34FA80";
    attribute INIT_3E of inst : label is "019B99B810305181F80A78E3463FA028C246BF3E80ABC80AB8FFA029D3C02529";
    attribute INIT_3F of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAF7F530F5FFF5FFF55FFF555FFF55";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "E288A09207DF0A2E2E22A82E0AAC82228BB028BCD3F08228840003001667F188";
    attribute INIT_01 of inst : label is "42A0A922FF888BA88888225998BFFFFFFFFFF42920AA2322E5B3E3E38A2E30F8";
    attribute INIT_02 of inst : label is "D22A6CFC6B82B86B82A823A208E8823A208E88BCF2AE2800B8BCF3A08208BCAC";
    attribute INIT_03 of inst : label is "20820820820820BBBBBBBB88888988888988AC186182082082EF3D00B4D34D34";
    attribute INIT_04 of inst : label is "2E61F08C2928A42A0A90888CCA0F367A098A8B2808888882220A86E088218608";
    attribute INIT_05 of inst : label is "184332393CD9E86838F0888ADA2B68691B8B8B899193CD9E8F92828A289890A8";
    attribute INIT_06 of inst : label is "09A83B2222616A2889898A49288A28890A82E5F083A1822F3EE23AEFCA22A682";
    attribute INIT_07 of inst : label is "322BE0AE200000FA50000000000000012927C3FF220A1A0A02223CB19FCC8FFA";
    attribute INIT_08 of inst : label is "C9F8CCC08CC082230A0000000007F8A288820822273BBFE993F8A22BE0AE8A22";
    attribute INIT_09 of inst : label is "2AA620AEA88CDC8CCC8C20A8708330B8F084223083E3CCE2A4C2924088BC2909";
    attribute INIT_0A of inst : label is "CA42290A88A888822331232230A808CCA5088230A8080B8B88C08C0830A86F3E";
    attribute INIT_0B of inst : label is "BCF09C363082B422376A022652E610B8B8AE089CC26B9888898DFA4C8ECE8CCD";
    attribute INIT_0C of inst : label is "FFF08822376F330822088A308C270AAEAB8330A8ACA48D9C22B98CDCDC2370A1";
    attribute INIT_0D of inst : label is "88DC8C2330A8330800550308A888E8ECCE10AF0BCCE30BCCC2B42208AD337233";
    attribute INIT_0E of inst : label is "308330A8F3CE13822CCCEA888EAC9E5F3CE23333AE82230DC270A123AB388220";
    attribute INIT_0F of inst : label is "F088FCCCEE232F30A92E3C8CBCC2B882238A08C230BCF088DC8DCAE3338BC222";
    attribute INIT_10 of inst : label is "0888888888888888888C888CC888CC8033014002D0888C20C2A932122842C20B";
    attribute INIT_11 of inst : label is "12A32A933F2392DA32302C8E4B68C8D54A8899886108C3308CCA82222222222A";
    attribute INIT_12 of inst : label is "F3C288BCFC6218862188A60E84C3BCF286889889AEE8B9898A800000000155E4";
    attribute INIT_13 of inst : label is "23EA0BB88233333622626F3C88188989BCF6F3DE898989422410408262622626";
    attribute INIT_14 of inst : label is "38BCFF8E28BA8A7CF0A22F7FCF55555522F3C60860899F3F3B8A2EF3FE820863";
    attribute INIT_15 of inst : label is "8FCF0888C2F1B9F9F9B3E822322723E272733EA0B82333330E30E2F3C28A988C";
    attribute INIT_16 of inst : label is "00055FA000000000FFAA550064E2E2E260E2E2E2F3C2222998A6625102302600";
    attribute INIT_17 of inst : label is "328720888A48A662438F9FCF0A608220888868966062823F30BF82E0A21A6E20";
    attribute INIT_18 of inst : label is "3FA4FEE0B82889EF3C2222E7BCF0888B9A4CFA0C8220A228720888A8B86E3323";
    attribute INIT_19 of inst : label is "000000000000050000422323B2BB3B2BAE08C88C2A0F8CEF8CCCEF8CCDCF8C27";
    attribute INIT_1A of inst : label is "CDCDCEB98249C8C8DCADF9932122B42C8620882AD5E2EFA88EBA22AAAAAAAA55";
    attribute INIT_1B of inst : label is "0AE26266F3F085226222000EB8220AE2E3C2108E2333882620F212212250B84D";
    attribute INIT_1C of inst : label is "46273AE0899883C848848842FC0BF022222002DA36FF39AE662336F3EE6B463B";
    attribute INIT_1D of inst : label is "0166BAC00000001DC0154008801928E6119CE3292B0AE62002938C27A4E237B0";
    attribute INIT_1E of inst : label is "2631A96708C262631A526708C2088C8BD822322F6626236666858260A4333380";
    attribute INIT_1F of inst : label is "BF30A8C2A408C2A408C2A40A0E2E2702702A4CCE30A9088C2088C20AE6727664";
    attribute INIT_20 of inst : label is "035410100004223B3324DC8A42290A20C08C08CE8830230233333AAA2A8882A0";
    attribute INIT_21 of inst : label is "2B829828829828828880000000000000143FA9503FA950121A884AA57895E420";
    attribute INIT_22 of inst : label is "9898F8E28B9CCAA3A22BE38888E189A2EF8E2899CCAA3A3E38A2A88B9FC6888C";
    attribute INIT_23 of inst : label is "401555555554015555AAAAAAAAAAA13F000000010FF588E3E38A2E6238F8E28B";
    attribute INIT_24 of inst : label is "55555596955569655969555696559556A9556559556C955655AA96A96AA55555";
    attribute INIT_25 of inst : label is "5515A9655556A550965A5960550965A596055A9555596A55555555555555556A";
    attribute INIT_26 of inst : label is "55955659556559556595565596955569655969555696555555A9555555555555";
    attribute INIT_27 of inst : label is "C61186D182221C20C61C8863FF3FF55555555555555555555555555AA96596AA";
    attribute INIT_28 of inst : label is "C604886B4221A86A0A82623083B42A09A208B87181221AD0886E1A82A0888C61";
    attribute INIT_29 of inst : label is "2F10C2882138BC2308E2085020B86E2F0B8622F08C2007CF08AA2B6220A82E21";
    attribute INIT_2A of inst : label is "82EB46888CC6E2BA5B8C618601186088CC231A20AA2F08E22F3FCCE28620882E";
    attribute INIT_2B of inst : label is "FCFCFCCFCCFCFCFCFED0A82E332233AE2BAB888F88EBFF23EF4621886E18220A";
    attribute INIT_2C of inst : label is "FFED960F281CAEAA3AA2AA22CA68A1AA0AA2CAABA3AA2AA22C8EB8AB8AC8B8FC";
    attribute INIT_2D of inst : label is "403FC00017C0003FFFBFC00017FFF400003FFFFFFFFFFFFC0000000000000003";
    attribute INIT_2E of inst : label is "C000002FFFC03FFD4001FFC000003FFD403FC00017C03FFD40003FC017FFC03D";
    attribute INIT_2F of inst : label is "00003FC0003FC000000CFF04000FF30001FFC03400003FC001FFC00034003FC1";
    attribute INIT_30 of inst : label is "05028500000528000000A0800020A00000002800000280000000050000050000";
    attribute INIT_31 of inst : label is "50003FC5003FC00005003FC0003FC0000028A0BC00E0A2B003CA280500428A10";
    attribute INIT_32 of inst : label is "00153FC1033FC001800FF00001400014000C2A40057E0B1500003FC5003FC001";
    attribute INIT_33 of inst : label is "40015C80003CA300000C92804173331550000BC000B8000000036FC1503FFC00";
    attribute INIT_34 of inst : label is "00A0002000A000000080000000941C141C003F005FFF003D40003F005FFF003D";
    attribute INIT_35 of inst : label is "60200BC0002C608000000BC0002C60000020002000A000000080000000800020";
    attribute INIT_36 of inst : label is "002555AAAA8000440554013FFFFFFFFC03C007FF00001541FD0000A000A02D5C";
    attribute INIT_37 of inst : label is "55F956FEAAF2AA3AAA8000054000002560115011101410104000000000000000";
    attribute INIT_38 of inst : label is "03C15505543FFFFAAAFBE0B820BFFC3800B8F03F0BF8FCB0BCBBFBFC00B5A5F1";
    attribute INIT_39 of inst : label is "003C03C007FF00001555557FFFD0003FFFC000400015557D0015557FFFD40000";
    attribute INIT_3A of inst : label is "8A228BFC68AE223D883B2E0EF3B2E138ECA2868ECA208A333288228CCF43BFBC";
    attribute INIT_3B of inst : label is "CE621A2889CE621A28888DCE621A28888CA62988610B3BA222A34A133390C3E3";
    attribute INIT_3C of inst : label is "08844054210015155484084150955400003AAAFFFFC820400000000155555555";
    attribute INIT_3D of inst : label is "0041500C440543304150CC4405433008468EA30C24CA020103A0415150C80015";
    attribute INIT_3E of inst : label is "0110110150055515015044044440054110540000150001500000054000154540";
    attribute INIT_3F of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEA0EFA0AAA0AAA00AAA000AAA00";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
