-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.Vcomponents.all;

entity VISIBLE_ROM is
  port (
    CLK  : in  std_logic;
    ENA  : in  std_logic;
    ADDR : in  std_logic_vector(12 downto 0);
    DATA : out std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VISIBLE_ROM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'    => result(i*4+3 downto i*4) := x"0";
        when '1'    => result(i*4+3 downto i*4) := x"1";
        when '2'    => result(i*4+3 downto i*4) := x"2";
        when '3'    => result(i*4+3 downto i*4) := x"3";
        when '4'    => result(i*4+3 downto i*4) := x"4";
        when '5'    => result(i*4+3 downto i*4) := x"5";
        when '6'    => result(i*4+3 downto i*4) := x"6";
        when '7'    => result(i*4+3 downto i*4) := x"7";
        when '8'    => result(i*4+3 downto i*4) := x"8";
        when '9'    => result(i*4+3 downto i*4) := x"9";
        when 'A'    => result(i*4+3 downto i*4) := x"A";
        when 'B'    => result(i*4+3 downto i*4) := x"B";
        when 'C'    => result(i*4+3 downto i*4) := x"C";
        when 'D'    => result(i*4+3 downto i*4) := x"D";
        when 'E'    => result(i*4+3 downto i*4) := x"E";
        when 'F'    => result(i*4+3 downto i*4) := x"F";
        when others => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO   : out std_logic_vector (1 downto 0);
      ADDR : in  std_logic_vector (12 downto 0);
      CLK  : in  std_logic;
      DI   : in  std_logic_vector (1 downto 0);
      EN   : in  std_logic;
      SSR  : in  std_logic;
      WE   : in  std_logic
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
    rom_addr              <= (others => '0');
    rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "9D031F8D0440640010402447C6464004308D900080530262C0C421153851B111";
    attribute INIT_01 of inst : label is "06B000EF62401449025540D46E6C000D000000002730340E360701101D09035C";
    attribute INIT_02 of inst : label is "C40B119B1009D324D4E25C62D3604B1EE134466EC1DA7B9119E4910CF511F7D4";
    attribute INIT_03 of inst : label is "13B8CF0B3244035C9D274CC92B3640358C91B407C50041C1C86B24C64040C309";
    attribute INIT_04 of inst : label is "000C000000000084000340000E00002C081D00D7000000919B1819013004191D";
    attribute INIT_05 of inst : label is "233302033223E102213FD032210087FDD83950282A773CB4003AC0005E000334";
    attribute INIT_06 of inst : label is "D9D3664C83A2B8A63E8A7EF3FC37EF3FFFFD00CBFFFC3FFFC64443FFFD323233";
    attribute INIT_07 of inst : label is "C47164301D27736BCF41B4035C9DD57334C2490D57306409243B017D05501DC4";
    attribute INIT_08 of inst : label is "400F70BE0D3C7CFF3C003CFF373CD589DB676DBB77579011111112026D800500";
    attribute INIT_09 of inst : label is "694134C414CD1818C0A450708BBB374A4641536A4C1DDD02C300A031AA274073";
    attribute INIT_0A of inst : label is "50C8614331C5230C86148C62A8042AC0AAA0036241416424A2DD1A3086265092";
    attribute INIT_0B of inst : label is "46222331C7186184858B47AA1117B49A0C011C41840099854754D4A21D51331C";
    attribute INIT_0C of inst : label is "4731C4731C54C40C91201DD1491277074200D8A1128C1D208CDD268244674447";
    attribute INIT_0D of inst : label is "AAA74535328C9070522A40232211DB5C575C4149C71D1C8C54C715881C71531C";
    attribute INIT_0E of inst : label is "249349A4080461C5D1011271011411859C4E031011C48904C68126408004D90D";
    attribute INIT_0F of inst : label is "07450C81D010D9D070B7908CB240241D1644070C03014D081104441D2234485D";
    attribute INIT_10 of inst : label is "630210810C226134164C206066AD12060CD833400A0145C041181C08341936A7";
    attribute INIT_11 of inst : label is "F10EB0E5B000024D3A41933E400013C43AC396C90601AF800080008A9E810C04";
    attribute INIT_12 of inst : label is "0008488E2BD4002006CE70080000D46DC006BC0C2447FCEF4050095B51AE4184";
    attribute INIT_13 of inst : label is "D900E106C71FFC08000300AFD100640EF35C3C08000000AF3D802880C856C020";
    attribute INIT_14 of inst : label is "4A1D7B135CD27638F35CB03E307691C37D71133C6844A8C6E4C3A80B8B4D400C";
    attribute INIT_15 of inst : label is "0864E94F46308A128F3647EB90D92942304F29A0DEB712B87B6E46C83512328A";
    attribute INIT_16 of inst : label is "E73B4C2362043B792439316DD38CC7924D1CB11E443F4C364FE102E238089152";
    attribute INIT_17 of inst : label is "A8CD91CC79E89E26E2466BD3939A6EE384B643324D1E0C90A5094D9CC7D64911";
    attribute INIT_18 of inst : label is "33661E394424389443909384341D338A50F949CD32031180F4FB9F1E4EF91349";
    attribute INIT_19 of inst : label is "00008844444000444888880000218311314388E74C8A4EDA0AB93A2435484398";
    attribute INIT_1A of inst : label is "4C00E40AC63216BF0A7C086F87A412F3653413E180002223921600D000000000";
    attribute INIT_1B of inst : label is "000000000000000000043930C708728914637806EA063182C444389340B03932";
    attribute INIT_1C of inst : label is "6A156012010868110E8990000406D902D85C1088141080D09981991251D11912";
    attribute INIT_1D of inst : label is "61D74E3615A69DB6695D0945351A476896615824568342914D4224892A748061";
    attribute INIT_1E of inst : label is "A2D1A918D15191DA1B8C55A5634065B495C511DD74E16DDA6D5D398907697144";
    attribute INIT_1F of inst : label is "D194AB5529B666130800C9B47DB76A5008A5125CD92115B7C964449D20980422";
    attribute INIT_20 of inst : label is "4449E33000BA94D811E69110340BA94D81502EA536066D5915F329DAA6800426";
    attribute INIT_21 of inst : label is "295510B4136249C623B374060B01D0A51110382449C024402354911766448B56";
    attribute INIT_22 of inst : label is "1715445C5410CF1070B01519D9005464290262580349112449D9098A5654454E";
    attribute INIT_23 of inst : label is "0B2CD1408D5150101981614851094148911076344DC9D813489912706449C151";
    attribute INIT_24 of inst : label is "924014B10602511D86811920264593641188C91730514140065586629821D442";
    attribute INIT_25 of inst : label is "36721716574642082430860475564474707658199591D5D991511D2158446411";
    attribute INIT_26 of inst : label is "68042855D0230D17648A99D055235DC18580F20A37744958596C95A8D4DDD328";
    attribute INIT_27 of inst : label is "D1D36355C115DD52D4705A6B4B51CD5169A69AD0DD85D0E0E4DD551E3881C241";
    attribute INIT_28 of inst : label is "1D772674950B0904D99923445D3606344D1453510348966A6740548D57061619";
    attribute INIT_29 of inst : label is "05D262AAAB766414113A4844574441411186055A175C1955DD5923447764815D";
    attribute INIT_2A of inst : label is "4299C87512448BB09DD1906B8D8BD1234DC941545115541C2452672A219809D1";
    attribute INIT_2B of inst : label is "706ABC24420A69B66A5CA61D876D99344944599461D24C21B71611B689535664";
    attribute INIT_2C of inst : label is "C41C1C0513498172C950475464744768800CC62998762916669D844824890204";
    attribute INIT_2D of inst : label is "E30315D66A74DCA095A05467745D9F6A47001DDDB2214A5412885152172C9DA3";
    attribute INIT_2E of inst : label is "85CB266CF148DC4941C230CA095A35A519DD24546470C04746CB04667647746C";
    attribute INIT_2F of inst : label is "2C1195D919D52AEB30411D9B2214A720D12E1505418853D82804487ACD148D14";
    attribute INIT_30 of inst : label is "C59151DD1C74755D2475374C50DDC88A8D9B28C5F10703077754677009115D1B";
    attribute INIT_31 of inst : label is "53D88044944AD02CC324454766C8D513230828DD19166A154D504A0C5B085526";
    attribute INIT_32 of inst : label is "A154901C5021411125140D5628DD254C35345180A374D2678D164DF6081DDD88";
    attribute INIT_33 of inst : label is "C1DD1955115D671D1F3448985F10700144DF40A081051700171607C41C005002";
    attribute INIT_34 of inst : label is "420635535818D54D601D6055DD60955098C498D0145F1070599151982114040A";
    attribute INIT_35 of inst : label is "15410811441451440428DD36A15450A01DB3051074D9094DD16374245462105F";
    attribute INIT_36 of inst : label is "5220A855240228DD172B448806314CCC0DD2C0D00840E0926A0700341D184404";
    attribute INIT_37 of inst : label is "88050C1837665515C83350C573154C5631400091A085D5050507540714D13007";
    attribute INIT_38 of inst : label is "0156AAFFFF0000000000FFFFAA9540F94FDBF8BFDDB00E4D571B00E77FE2FE7F";
    attribute INIT_39 of inst : label is "000000000000101111110000000000000000000000000011100332211000016F";
    attribute INIT_3A of inst : label is "FFFFFFFA4E4E794888B72CB1B1BC5ABF0000003FEA513E943001111111111110";
    attribute INIT_3B of inst : label is "FFAA50E70D1E4E53A53E94016BC45A8FC000000CEA53E4E4E38DE22216DB1B1A";
    attribute INIT_3C of inst : label is "394E5393E4E4393EAA955400FFA9543EA50F94F93939E340000000100000000F";
    attribute INIT_3D of inst : label is "254C03FFFFFC1CA53C34CBF4F93F0006206201B400021050FA50F943E53E53E4";
    attribute INIT_3E of inst : label is "06418D990A4709118E5000940D980679719100911CFFF377624DA80D14020265";
    attribute INIT_3F of inst : label is "DB35F214F022010C08A8851511A222AAAAAAA95557FFFFD55005A80AAAAA8C40";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "1E00C310301173001040054F0817300410024002AA0FF83011860B2E38F30022";
    attribute INIT_01 of inst : label is "1830003FCB40211D001AC0190D070012700000003434490C43270690141C1994";
    attribute INIT_02 of inst : label is "06472641190D003819C35543E4050710D0089905810446F4305CF40D3B1004EC";
    attribute INIT_03 of inst : label is "2DF1078F074519941E3400DE1707B19810E17C77499185E64D83381730641F8D";
    attribute INIT_04 of inst : label is "000680001900001000008000050000100C140665000000E641205CC03476101E";
    attribute INIT_05 of inst : label is "100011230133C133003FE022222247CB6B330231ED2FAFC40015000064000090";
    attribute INIT_06 of inst : label is "D5C3560E609375E5B1FC3D3FF242DA7FFFFC2133FFFF3FFFF01303FFFC331101";
    attribute INIT_07 of inst : label is "8039EC301407B44300713C19941EFB2008D05D0FB2017301742E1954659D9A80";
    attribute INIT_08 of inst : label is "000FA3FFCCFF3ED7BF00FCFF3382CD023C5F0000070392E2223332143400003A";
    attribute INIT_09 of inst : label is "C772A68CD009A0E49CAC806376661A684A5794E963DA9E7D0A1795C247059761";
    attribute INIT_0A of inst : label is "95F8A257E289501F8A25806EA404EAC0AAA04880920146DAAA128030040958DF";
    attribute INIT_0B of inst : label is "4A129122AA28AA8A57A4A56AE96D55350C8B28B2880887444776DCD81D127E28";
    attribute INIT_0C of inst : label is "89023880238A380C56989A5205695629692244A932A49AA44545F9415A694948";
    attribute INIT_0D of inst : label is "AAA5A2B90B80D282A6160CA9202778B288B1A60A18A924018A18220061862860";
    attribute INIT_0E of inst : label is "3DB3D79444A20A4999426A5228289A49E4098122824C55C01D6A6232900A6989";
    attribute INIT_0F of inst : label is "2D96088B602C25819238A8C2CB88B22D2B5A28B2F122B2CC934E0C3EA2DCA07E";
    attribute INIT_10 of inst : label is "AA00D242C4928209095F7C81956BC1093021C390407146C0C328ED0C35FD6E95";
    attribute INIT_11 of inst : label is "522D7875DC0003FB3DD77EE500001C346090820208F60FC000C000CFC5CDC837";
    attribute INIT_12 of inst : label is "0001078283C00040052187F3000026E2C0181C00054F403FC084006464162888";
    attribute INIT_13 of inst : label is "C0003001411103F30001A362C400B800054143F3000191603C001D0066001FCC";
    attribute INIT_14 of inst : label is "9920E44210801438C338B93FD2B6F9030EC242A44F629527A5059105818684E4";
    attribute INIT_15 of inst : label is "B8D53A128FFE123DF8148EA402523A5493913810E55301C4E3D55300943D2953";
    attribute INIT_16 of inst : label is "554290099CE4143E93951690F3C669540F25DE90CA4DA3280DFF4F53EB3F63D2";
    attribute INIT_17 of inst : label is "52D000753D0C4574F15174F1540750F325DBC397FAA30E57AA00A68C0A580542";
    attribute INIT_18 of inst : label is "4397C03CA5C035F30954FC3015C31687C06CA506170195C07F814F0553C0015C";
    attribute INIT_19 of inst : label is "DFDFFDFDDFDDFDFDFDFFDF0000E384E2935D4FAE534EFA54CEEA94D53BA753E3";
    attribute INIT_1A of inst : label is "0F2FFF07C040F70013EB643A156A0FB017EA3EFFFC0011115515626000000000";
    attribute INIT_1B of inst : label is "00000000000000000008EA98BD8FD1CE80FEE8000000300BCF0AD4AD53A5402C";
    attribute INIT_1C of inst : label is "1EC4B72B72849899A9099A0A40A0B8C8B0E424502C2454E0C50AD52A96929920";
    attribute INIT_1D of inst : label is "4F1FA024F93C393E4F920262B9178FBC3E4F9E38EBC08098AE45244121E40F77";
    attribute INIT_1E of inst : label is "A07A07289692996EC73016184390463E84C12191FA024390C31FE44606433048";
    attribute INIT_1F of inst : label is "B80E02C9072D832F4CA4482E372DAA280083284C1A41211FF0E6666C030CF092";
    attribute INIT_20 of inst : label is "6666D334002D0AE82D9999A02402D0AE82900B42BA0A4B2996FC0721C30C04A0";
    attribute INIT_21 of inst : label is "899D2248EBA380F1185078414A20E041A1220706A1488002A38731CC784802CA";
    attribute INIT_22 of inst : label is "A52A6694A5070E10B450999555A15562C521184790611C048DDD8B76766769C9";
    attribute INIT_23 of inst : label is "8D14922C892924949ACA41A4EDCE71A4ADB3A42A698A909A68A99A52A6694A99";
    attribute INIT_24 of inst : label is "6A408A220A00D2D28DCDD6833E87E3F89E2F0A890050000014750E406A02113C";
    attribute INIT_25 of inst : label is "06804A04484A3C8C00108434A7B6B4A4923BAC9A999292DEDAD6D22CAB08DCDD";
    attribute INIT_26 of inst : label is "640A2692E830B227642999E852127E1DDC4A2C410486C1241618161410112805";
    attribute INIT_27 of inst : label is "53A98184C12191932130461A4C84C1911861869091491C1010919123C0420C42";
    attribute INIT_28 of inst : label is "99F976489D80311B5959127772860B1842362B902564366667A14849E8777199";
    attribute INIT_29 of inst : label is "BADE955555595624291555795495624291560844084C1919195D136766644D9D";
    attribute INIT_2A of inst : label is "90618084624848620E121883028B72838E08635ADD375AD0C463322A91540D55";
    attribute INIT_2B of inst : label is "90AAAB2480290B1D2A102CB53B4A5595A860522C8BE044A41C14E52AA8724976";
    attribute INIT_2C of inst : label is "882D2B4A1383A2B10D235A64A494A79B0AEB01061085210584610844943C07E4";
    attribute INIT_2D of inst : label is "5D00310C686418181650844768D5D1C44AC09E5E411281E82044A03A2B10D26F";
    attribute INIT_2E of inst : label is "8AC434974E84E2C282B3108141650B1111DA35B644AC4259490A0485B4A49490";
    attribute INIT_2F of inst : label is "28121AD29252AA942C4925E411283E28A9292A0A824CA3F4DA2A48A504E84E2E";
    attribute INIT_30 of inst : label is "0111292520F483190486392914E4845549641B02E20B49E4949497ACC9969524";
    attribute INIT_31 of inst : label is "A3FCA2A494A5B110B0265A494908E129D72390559715A4266688A92010C0A13A";
    attribute INIT_32 of inst : label is "4266602488DA2D28190806DDD0999AF0A112D20A415663EB021C8F1B67925244";
    attribute INIT_33 of inst : label is "89252929A120E83D24E4ACA02E20B41284E2C0231E792823182A0B882D0A8482";
    attribute INIT_34 of inst : label is "823B03D838EC0F60D790EFD250E392932C80982CE0EE20B4DA92932C11284F02";
    attribute INIT_35 of inst : label is "A2220C1204A0A208049055B64266681C2DB02829641A418E48439025A4B11280";
    attribute INIT_36 of inst : label is "E0029099988090558706C00545A28941CE4A91B14060BD521196F90659C14844";
    attribute INIT_37 of inst : label is "2205206C37B79715B4C08B0E0C38F020C088DA821783E283C20F8A0E38B11284";
    attribute INIT_38 of inst : label is "AAAAAAAAAAFFFFFFFFFFAAAAAAAAAA555FF939DDD861BC6B0E93E4927776C6FF";
    attribute INIT_39 of inst : label is "1999111911918008088000808080808080808080808080833332222222208555";
    attribute INIT_3A of inst : label is "FFFFFFFFFAA540FA50E94F94E93A4E4E9393938E4E4E79393199119191919191";
    attribute INIT_3B of inst : label is "55555503EF34E3924E793906C6DB1B2B2C6C6C681B1AC6B16F16B05AF015AAFF";
    attribute INIT_3C of inst : label is "955003FEAA55403FFFFFFFFFAAAAAA95555000FFEA9503C00000002AAAAAAAA5";
    attribute INIT_3D of inst : label is "666406AAAAA35A9FEBE52AAA4548000050050400B48B78FFAAAA5554003FFEAA";
    attribute INIT_3E of inst : label is "0751C1C10C5001618030090401D40841F5CE00153F6AAFE65F710001EC020242";
    attribute INIT_3F of inst : label is "D37FC0A000F08B2C3C29F1159255551555550005400055400555555555554D70";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "51000054A109004038E291502510068E2BE068A2AA5B0442AA69806FB2C80CA8";
    attribute INIT_01 of inst : label is "904AAA40122A9008A9042A501D12801428000000058650015293044000809006";
    attribute INIT_02 of inst : label is "6060944481080582400005080415008108925110A8015284844A849160841182";
    attribute INIT_03 of inst : label is "9005640090109006512016108090010056084204441925046904025006064001";
    attribute INIT_04 of inst : label is "FFFFEBFFFFAFFFFEBFFFEAFFFFABFFFEA680A401AAAA8A944412401886000491";
    attribute INIT_05 of inst : label is "000000001113C000003FD100011043E9CA622121DE5B3323FFFFEFFFFFBFFFFE";
    attribute INIT_06 of inst : label is "000000000184310005403FFFFC02C03FFFFC0023FFFF3FFFF31233FFFC001200";
    attribute INIT_07 of inst : label is "0034ABFA80947414250840100651DEDA8119100DEDA90064403B0C0120008000";
    attribute INIT_08 of inst : label is "E6400341CCFF3F00FDEB7CFF33FFC00882007FB5B7579226AE2222000000003F";
    attribute INIT_09 of inst : label is "E9339B7749B4E3C34E0B72A99999F1AA092749E1A44E4EA2A9A4690DA8E0A8AA";
    attribute INIT_0A of inst : label is "6A0451A811469C20451A7080032800720007288485CA29CE06928850A8C1A24F";
    attribute INIT_0B of inst : label is "08E40C1545155145AB9099A0E4AD9236294114D14CA92922A919614284828114";
    attribute INIT_0C of inst : label is "495144B554494CA982634642182690D195405908E42346075A78FE8A09190A0A";
    attribute INIT_0D of inst : label is "80119270D3F4CD0D19D83D00CC13F9644944FE544D1427144B4D1253C4D12534";
    attribute INIT_0E of inst : label is "42F42F92FD264328B87C2EF7C9238E386294AF7C92296A215591A2340C0A26D6";
    attribute INIT_0F of inst : label is "4563E3D15E2306E8B476F65514D026282E0B2D652B4267A991454516B4748902";
    attribute INIT_10 of inst : label is "A7E24AE663B8A84141A8B08419AC14D3010D041F8B4C109410210EA8A2789E1B";
    attribute INIT_11 of inst : label is "857A05E812AAA957FFA07FFFEAAABA05E817A05E813411AAAAAAAAAA91A4AF92";
    attribute INIT_12 of inst : label is "FFFFE6A1ABFEAAFAAFFFFAAFAFFFF1A1EA904292915003402A42A41D4063E15F";
    attribute INIT_13 of inst : label is "FFAAEFAFFFFFCAAFBFFFF962FFAAEEA3FFFFCABEBFFFFA62BFEABBEAFFFF2ABE";
    attribute INIT_14 of inst : label is "38290FFE00943FE80EE8803AA1A4EAA18A543E90A0E4CFD40004D544C4C3C0F0";
    attribute INIT_15 of inst : label is "807FEAE8042AE813ABEA04AFFEA812FA013813C3403E2B30A803FE093FE82BA8";
    attribute INIT_16 of inst : label is "AAA9551AE2552543A95517AA54097AAAA01532AA0553A81553A284FEA810E13E";
    attribute INIT_17 of inst : label is "A30053800050B00103FE0103FFF88500FA0404F8001413A81445F9505DA54557";
    attribute INIT_18 of inst : label is "02A80020AA00EA000AAB0000EA00283003800008C00E03038003C03800001003";
    attribute INIT_19 of inst : label is "7665647776666766565774000000000002000AA0000A00000A00000028000220";
    attribute INIT_1A of inst : label is "0F10FF16BFF1A6FF140AD442FD5512AFFEA52A02A80011113D30D15000000000";
    attribute INIT_1B of inst : label is "000000000000000000000000000000003C00000FCF3C2C028A00800800000300";
    attribute INIT_1C of inst : label is "EA30A02E0EE9A98A5A18A51A12A5E919C70F01470FC143C2B410A42886868822";
    attribute INIT_1D of inst : label is "1E0DEDA1E4790A719C6E8A9270FA2DEE719C69A2FEEBA2A49C3EBBEDA4F24F3B";
    attribute INIT_1E of inst : label is "0D149422464644EA3A81C244878C917A3B6020A0DED9128490282080CA12D808";
    attribute INIT_1F of inst : label is "E55C2708537092C2A92305797F70A024AD15E4B60220204EC491196A90434D34";
    attribute INIT_20 of inst : label is "1196BBAABE7089C10A66442FABE7089C10AF9C2270429C2442B0D425924AD295";
    attribute INIT_21 of inst : label is "2CCC2BBA27850B82240C3ADA3349E2286829595096D015CA9F13B4ED1908A709";
    attribute INIT_22 of inst : label is "E85229A14FBC3D8C3ACA0220225800AE08C22C3C44B2D180ACCE93B33BB39E1C";
    attribute INIT_23 of inst : label is "ABB202F3E02821838210E8B34A18E8934A462042BA1483A69148AE85229A148A";
    attribute INIT_24 of inst : label is "66D409C9C022868E161466784390240AD0B036484AC00000B3BCEC051051EED3";
    attribute INIT_25 of inst : label is "719F8B730B0AD3A8B2CBEC9090A1A0A1B477B6828802028E82464E852A61A18A";
    attribute INIT_26 of inst : label is "13C05242C5470EA9389ECCE1C2FB37ECEFAAF32EB0BB5C27C2E9C2E5E9CE2678";
    attribute INIT_27 of inst : label is "4BBA860B6020A06BB2D80822ADCB6060208208AD803623070F80602F36F0F3E9";
    attribute INIT_28 of inst : label is "6CDDB1BAA64BCFB8868EFB1B37A1C1D3AEA9270C19B093BB33870BECFFB3BE46";
    attribute INIT_29 of inst : label is "734CEA22220A2BE1E4EAA23AA0A2BA1A46A2E088D2B60E0E0A8EFB3B1B3BEC6C";
    attribute INIT_2A of inst : label is "B51ED47BBC0AD2B49E86888B66D1D22BAE339A0BA8A2898F3EE95F4ACEBE24AA";
    attribute INIT_2B of inst : label is "852ABC80BF425E56E0E271F865998A68A3A3A2739C22DF095CA1B86E239C0A1B";
    attribute INIT_2C of inst : label is "6F0EB0DD8F2FA2CB28291910919393B429201E91E47B4FB0B13C4ED0364CAB20";
    attribute INIT_2D of inst : label is "E3299E67A0B2C52702E9B2B1BA4A4AC80BE2CECECB5B6AF622DEDAFA2CB282D3";
    attribute INIT_2E of inst : label is "8B2CA0BCE363CBCB62F8B252302EA32CAC6E909280BE2B1B0B2CB080A0B1B2B2";
    attribute INIT_2F of inst : label is "B2C20286CACA40ACBE6CAC2CB536BCAD24CA2D8B62D0DBF2CB4930AB2C363C9E";
    attribute INIT_30 of inst : label is "68EC2C6CE7209CECB0B2F0CACFC330AA982CB430DBC3AF0280A0A3BE6CC6CC2C";
    attribute INIT_31 of inst : label is "DBF2B49320AAE8B2FAB31B0B0B25E82F23B0210269E0B87392D393638F08B4AB";
    attribute INIT_32 of inst : label is "8519650D5781C8ADF16294AA61465BC3159E82D18519640B6640909EB80A02D4";
    attribute INIT_33 of inst : label is "2C6CE464EC2709C82F23BBCDCDBC3AB763C9C8B4D3082FA4C1D0D36F0EA85189";
    attribute INIT_34 of inst : label is "CB8E9CEDEE3A7397B087BCC287B882F8B657A90F0F0DBC3AC282FAB6B4B64C8B";
    attribute INIT_35 of inst : label is "37D223C2D0368778ADE1CE6B873927070ADB4DE7B2C22C7CF32F3CB1B0AF40DB";
    attribute INIT_36 of inst : label is "B2B461465A32E1CE48C3A21210676E32BCF8C2E88A8AC38CEEF3447BED1B0AD0";
    attribute INIT_37 of inst : label is "F2E4A228A3A290D3CC043014D053C14F052D6A82FC9062521440894852EB4A06";
    attribute INIT_38 of inst : label is "000000000000000000000000000000000FFFEA50FA4390E401B06C1AF05ABFFF";
    attribute INIT_39 of inst : label is "88C4C800040844C0084C8400CC884400CC884400CC8844011111111111110000";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFAAAA555000FFEAA55003FEA9500FFA954030C80800CC884400";
    attribute INIT_3B of inst : label is "555555540E2A5403FA954000156AFF0056ABFC0155AABFF000555AAAAFFFFFFF";
    attribute INIT_3C of inst : label is "55555400000000000000000000000000000000FFFFFFFE800000001555555555";
    attribute INIT_3D of inst : label is "555007FFFFFBAAAABFAAABFAAAAC0000040040000B4940AAAAAAAAAAAA955555";
    attribute INIT_3E of inst : label is "0054050501510445050001400504054434020045421FFEEBAEA0000400FFFFE1";
    attribute INIT_3F of inst : label is "C4000BFE0902DB4E42AACCC48200000000000000000000000000000000000144";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "03000001000000C01862AAAAEAAAAE861AAFD8659982D4AAE34C0A2F38E3F188";
    attribute INIT_01 of inst : label is "AABAAAAAEAEAABABAAAEAAAABC05000050000000010001000D0F003000000000";
    attribute INIT_02 of inst : label is "4000000001000000000000000000000000000007AAAABEABAAFAABABAAAAAEAA";
    attribute INIT_03 of inst : label is "0000000000000000010000000000000000000000000000004000000000000000";
    attribute INIT_04 of inst : label is "000000000000000000000000000000000EAAAAAAAAAA80000000000000000000";
    attribute INIT_05 of inst : label is "000000000003C000003FE000000323CF43213130338812300000000000000000";
    attribute INIT_06 of inst : label is "000000000000140000003C17D001403FFFFC1213FFFC3FFFD11033FFFC000000";
    attribute INIT_07 of inst : label is "4037003000007000C0300C000001C0000000010C000000000404000000000000";
    attribute INIT_08 of inst : label is "4AA00B3CECFF3C003CFF3E3CB07D000000010000032B92AEA662220000000005";
    attribute INIT_09 of inst : label is "88A28CAB3AB35232324B22A0CCCFDCA888A228A1A1222EA6492D3B4CCCCDA9A2";
    attribute INIT_0A of inst : label is "4A90812A42008CE90802339703B975330002388C808884AA5A00888C8A8DA828";
    attribute INIT_0B of inst : label is "8BFFCDCA18228609A29819E5C6899A662FFC2082089FC008488422122222A420";
    attribute INIT_0C of inst : label is "88C3088C3084089B22333222F21088FC4B9F2F04FD53327323228888888888A8";
    attribute INIT_0D of inst : label is "85594134C23088D9D9D83F9C8CDA68208820CA2708262F308C082222B0821020";
    attribute INIT_0E of inst : label is "8A68A699FC882A22223B30B3E2223A3322B6F33E222F69520DAD883E4CEA0636";
    attribute INIT_0F of inst : label is "E3A623F8E22336B0BE3AE2F0C3F3DA26098C08208BE0AE2FE28A0822BF388A2E";
    attribute INIT_10 of inst : label is "AA8266422390888C8DA9948CD9FA4CDE537A4DCDCA963BF8A1A3BF181A268A1B";
    attribute INIT_11 of inst : label is "5515545552AAA957D55555FFEAAA955455515545550AA8AAAAAAAAAAB0C61A18";
    attribute INIT_12 of inst : label is "AAAAA0A063CAAAAAAA8AA000AAAAA020EAAA8AA2AAAA20AAAAAAAAA2AA815545";
    attribute INIT_13 of inst : label is "CAAAAAAAA8AA8000AAAAA820CAAAAAA2A8AA8000AAAAA820BCAAAAAAA8AA0002";
    attribute INIT_14 of inst : label is "C03FF50000FFD500F040FFE403DF8003C7FFD400FF70B540000F800F8F8E0FAC";
    attribute INIT_15 of inst : label is "80EAAA000FEA003EA8000FA000003E0003C03D03FF103DC0FFCD000FD4003DFF";
    attribute INIT_16 of inst : label is "A900003AA4003FFEA0003EA0000FEA80003FEE800FFEA03FFEA20FAAA83CA3EA";
    attribute INIT_17 of inst : label is "A95502AA9500AA9402AA9402AAA99003AA500FA955403EA9410FA800F8A00FFE";
    attribute INIT_18 of inst : label is "52AA652AAA54AAA94AAAAA94AA992AA952A5AA8AA94AA952AAA9542AA95542A6";
    attribute INIT_19 of inst : label is "33331033210012333110000000514A5152A54AAAA94AAAA64AAAAA552AA952A9";
    attribute INIT_1A of inst : label is "5015001555015555155540555000155540000055540000004005000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000455545545514540555405451414054505545551555415";
    attribute INIT_1C of inst : label is "2A48A5725B1B7A658726583E32D826FC22327332B2F337F2623F622A6A626622";
    attribute INIT_1D of inst : label is "8268AA08220862088229084134CA88A408822A289A4642104D324AC8208908AA";
    attribute INIT_1E of inst : label is "CC7886226A62662A4E5332198F8D860A0A0626268AA0862186684554D8868189";
    attribute INIT_1F of inst : label is "261B2088C6088686CFF33609A208A0109CC6D1A06226261A9199942A061A1FF3";
    attribute INIT_20 of inst : label is "9942B3A8640884D2B27766E90A40884D2B29022134AC82266694C721C619F3D8";
    attribute INIT_21 of inst : label is "222224E4D10ACA155149D9F73FF6E2262627DF9846F3D98BCFDAA6A989889089";
    attribute INIT_22 of inst : label is "08FC84237B2D3B0CFC81656656C595B850E441A101C6B4989212FC0084884221";
    attribute INIT_23 of inst : label is "C92062B686222323323780C3F2338043720CC88CC23F22108372308FC8423723";
    attribute INIT_24 of inst : label is "22F3C4A0FE22626A3726522588A2E8A9A4A92108CD2000004A22898C38C32296";
    attribute INIT_25 of inst : label is "CD8C08C8888B96C824A2890B89898889BE3AA2222262626A6E6A6A66299F7E65";
    attribute INIT_26 of inst : label is "8BACCB21D0869904888321E332B0A222A895860248C8F223323F3233232120CC";
    attribute INIT_27 of inst : label is "26E888DA0626262666819554989A062655555522362162424236262B68F386C4";
    attribute INIT_28 of inst : label is "228888A4120A1B252222B088AE88CC8EC904134CC888888C878CCAC2988AA222";
    attribute INIT_29 of inst : label is "2A6A880444808C2310C880B08808C2310C8A8D9C8CA062626222B088888AC222";
    attribute INIT_2A of inst : label is "9C3270C8BDC9FDFF6E62688BCAFCE2269624848C224848286C9193F50CA02611";
    attribute INIT_2B of inst : label is "8DFFE958BF2D8209A022082609826500A0B3020B8222CFB60898260A208DC993";
    attribute INIT_2C of inst : label is "CF3F29F90FE2A2824224A88888898AA519653742208BFB08882209F3E0089948";
    attribute INIT_2D of inst : label is "8604E238A1A02F7372B08888A02229998A422A2293CE48A422FF922A28242296";
    attribute INIT_2E of inst : label is "8A0908A59643FB8A4290A0F7372B26622228088898A424888A4A089888888BA4";
    attribute INIT_2F of inst : label is "282262222A290B292422A2E93CE488AF10F2290A42F392222BC43C8A4A643FAA";
    attribute INIT_30 of inst : label is "82222222E3888E280889FDA227F6F323E3292537B3CFC85A99888BA422222229";
    attribute INIT_31 of inst : label is "9222BC43C8B290A4908888888A4BE2284BA572650CCC8C88422E4BF2384888AA";
    attribute INIT_32 of inst : label is "C884233F233CA2709C9DF32332210A10888A22F8C884288BCA8BA2A8A16A66F3";
    attribute INIT_33 of inst : label is "8222E222A22388E22948CE3E3B3CFC7E43FA88A1A6D22A3CDCDCDECF3F1F23C8";
    attribute INIT_34 of inst : label is "8A1B0E30E86C3843A923A12223A122A1AC332F73737B3CFC2222A0AC7CE4088A";
    attribute INIT_35 of inst : label is "C84A2332F3C88CC89B322108C884237332B32210A02222FF2CBFC888888FCF2B";
    attribute INIT_36 of inst : label is "627E322109F2322118DE4236253E42373F2A269189A1840F000A100C284889F3";
    attribute INIT_37 of inst : label is "F1D260281A9B88CED94DE93BA4CE53B94CDF7F22E1E20122338A0488CD83CFDA";
    attribute INIT_38 of inst : label is "000000000000000000000000000000000FFFFFFFAAA95500000556AAAFFFFFFF";
    attribute INIT_39 of inst : label is "666262A66A2AA6E6666EEEEEAAAAAAAA66666666222222208080808080824000";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAA955555550000000322226EEAAAAAAAA";
    attribute INIT_3B of inst : label is "55555555501555540000000000000055555556AAAAAAAAAFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "0000000000000015555555555555555555555500000000000000001555555555";
    attribute INIT_3D of inst : label is "3333F3FFFFFFFFFFFFFFFFFFFFFC000000000000400400000000000000000000";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFF157FFFFFFFFF0";
    attribute INIT_3F of inst : label is "EAAAAAAA8622FFEE8BBE56622200000000000000000000000000000000003FFF";
  begin
    inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
